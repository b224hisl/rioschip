magic
tech sky130B
magscale 1 2
timestamp 1662997953
<< viali >>
rect 101689 27625 101723 27659
rect 9689 27557 9723 27591
rect 10517 27557 10551 27591
rect 19257 27557 19291 27591
rect 22661 27557 22695 27591
rect 39129 27557 39163 27591
rect 43177 27557 43211 27591
rect 43913 27557 43947 27591
rect 45017 27557 45051 27591
rect 53481 27557 53515 27591
rect 61853 27557 61887 27591
rect 69397 27557 69431 27591
rect 74641 27557 74675 27591
rect 81265 27557 81299 27591
rect 81817 27557 81851 27591
rect 82553 27557 82587 27591
rect 86233 27557 86267 27591
rect 87061 27557 87095 27591
rect 87705 27557 87739 27591
rect 96537 27557 96571 27591
rect 97181 27557 97215 27591
rect 98009 27557 98043 27591
rect 100401 27557 100435 27591
rect 102517 27557 102551 27591
rect 103161 27557 103195 27591
rect 106105 27557 106139 27591
rect 108313 27557 108347 27591
rect 109417 27557 109451 27591
rect 110889 27557 110923 27591
rect 113649 27557 113683 27591
rect 115581 27557 115615 27591
rect 2421 27489 2455 27523
rect 4997 27489 5031 27523
rect 6377 27489 6411 27523
rect 7573 27489 7607 27523
rect 8125 27489 8159 27523
rect 30757 27489 30791 27523
rect 33333 27489 33367 27523
rect 34713 27489 34747 27523
rect 40417 27489 40451 27523
rect 41705 27489 41739 27523
rect 49341 27489 49375 27523
rect 54309 27489 54343 27523
rect 54493 27489 54527 27523
rect 63233 27489 63267 27523
rect 68753 27489 68787 27523
rect 71329 27489 71363 27523
rect 75193 27489 75227 27523
rect 79149 27489 79183 27523
rect 79333 27489 79367 27523
rect 85037 27489 85071 27523
rect 90649 27489 90683 27523
rect 94881 27489 94915 27523
rect 99113 27489 99147 27523
rect 107485 27489 107519 27523
rect 107761 27489 107795 27523
rect 108129 27489 108163 27523
rect 1593 27421 1627 27455
rect 2697 27421 2731 27455
rect 4261 27421 4295 27455
rect 5273 27421 5307 27455
rect 6653 27421 6687 27455
rect 7941 27421 7975 27455
rect 11621 27421 11655 27455
rect 12449 27421 12483 27455
rect 14289 27421 14323 27455
rect 15301 27421 15335 27455
rect 15577 27421 15611 27455
rect 17233 27421 17267 27455
rect 17877 27421 17911 27455
rect 19441 27421 19475 27455
rect 20177 27421 20211 27455
rect 20361 27421 20395 27455
rect 21005 27421 21039 27455
rect 22201 27421 22235 27455
rect 22845 27421 22879 27455
rect 23857 27421 23891 27455
rect 24593 27421 24627 27455
rect 25329 27421 25363 27455
rect 26985 27421 27019 27455
rect 28089 27421 28123 27455
rect 28825 27421 28859 27455
rect 30481 27421 30515 27455
rect 31401 27421 31435 27455
rect 32597 27421 32631 27455
rect 33609 27421 33643 27455
rect 34989 27421 35023 27455
rect 35909 27421 35943 27455
rect 36461 27421 36495 27455
rect 37749 27421 37783 27455
rect 38669 27421 38703 27455
rect 39313 27421 39347 27455
rect 41521 27421 41555 27455
rect 42441 27421 42475 27455
rect 43361 27421 43395 27455
rect 44097 27421 44131 27455
rect 45201 27421 45235 27455
rect 47041 27421 47075 27455
rect 48145 27421 48179 27455
rect 50537 27421 50571 27455
rect 51181 27421 51215 27455
rect 52201 27417 52235 27451
rect 57161 27421 57195 27455
rect 58357 27421 58391 27455
rect 58633 27421 58667 27455
rect 59829 27421 59863 27455
rect 60565 27421 60599 27455
rect 60841 27421 60875 27455
rect 62037 27421 62071 27455
rect 63509 27421 63543 27455
rect 64705 27421 64739 27455
rect 65809 27421 65843 27455
rect 66453 27421 66487 27455
rect 67097 27421 67131 27455
rect 67833 27421 67867 27455
rect 68661 27421 68695 27455
rect 69305 27421 69339 27455
rect 69581 27421 69615 27455
rect 70225 27421 70259 27455
rect 71973 27421 72007 27455
rect 72249 27421 72283 27455
rect 76113 27421 76147 27455
rect 76757 27421 76791 27455
rect 77033 27421 77067 27455
rect 80069 27421 80103 27455
rect 81081 27421 81115 27455
rect 82001 27421 82035 27455
rect 82737 27421 82771 27455
rect 83841 27421 83875 27455
rect 86417 27421 86451 27455
rect 87245 27421 87279 27455
rect 87889 27421 87923 27455
rect 88993 27421 89027 27455
rect 90557 27421 90591 27455
rect 91845 27421 91879 27455
rect 95709 27421 95743 27455
rect 96721 27421 96755 27455
rect 97365 27421 97399 27455
rect 98193 27421 98227 27455
rect 99389 27421 99423 27455
rect 100585 27421 100619 27455
rect 101873 27421 101907 27455
rect 102701 27421 102735 27455
rect 103345 27421 103379 27455
rect 105369 27421 105403 27455
rect 106289 27421 106323 27455
rect 107301 27421 107335 27455
rect 108497 27421 108531 27455
rect 109601 27421 109635 27455
rect 110245 27421 110279 27455
rect 111073 27421 111107 27455
rect 112453 27421 112487 27455
rect 114753 27421 114787 27455
rect 116041 27421 116075 27455
rect 117329 27421 117363 27455
rect 117605 27421 117639 27455
rect 4445 27353 4479 27387
rect 9413 27353 9447 27387
rect 10333 27353 10367 27387
rect 11161 27353 11195 27387
rect 11805 27353 11839 27387
rect 12173 27353 12207 27387
rect 32781 27353 32815 27387
rect 36277 27353 36311 27387
rect 36737 27353 36771 27387
rect 37933 27353 37967 27387
rect 40233 27353 40267 27387
rect 46029 27353 46063 27387
rect 54217 27353 54251 27387
rect 54953 27353 54987 27387
rect 84853 27353 84887 27387
rect 84945 27353 84979 27387
rect 89361 27353 89395 27387
rect 92765 27353 92799 27387
rect 94789 27353 94823 27387
rect 104725 27353 104759 27387
rect 1409 27285 1443 27319
rect 12541 27285 12575 27319
rect 14105 27285 14139 27319
rect 17325 27285 17359 27319
rect 18107 27285 18141 27319
rect 20821 27285 20855 27319
rect 22017 27285 22051 27319
rect 23673 27285 23707 27319
rect 24409 27285 24443 27319
rect 24961 27285 24995 27319
rect 25421 27285 25455 27319
rect 25881 27285 25915 27319
rect 27169 27285 27203 27319
rect 27905 27285 27939 27319
rect 28457 27285 28491 27319
rect 28917 27285 28951 27319
rect 30113 27285 30147 27319
rect 30573 27285 30607 27319
rect 31493 27285 31527 27319
rect 38485 27285 38519 27319
rect 39865 27285 39899 27319
rect 40325 27285 40359 27319
rect 40877 27285 40911 27319
rect 41153 27285 41187 27319
rect 41613 27285 41647 27319
rect 42625 27285 42659 27319
rect 46121 27285 46155 27319
rect 46857 27285 46891 27319
rect 48237 27285 48271 27319
rect 48789 27285 48823 27319
rect 49157 27285 49191 27319
rect 49249 27285 49283 27319
rect 50353 27285 50387 27319
rect 50997 27285 51031 27319
rect 52009 27285 52043 27319
rect 53205 27285 53239 27319
rect 53849 27285 53883 27319
rect 55505 27285 55539 27319
rect 56425 27285 56459 27319
rect 57253 27285 57287 27319
rect 59645 27285 59679 27319
rect 64521 27285 64555 27319
rect 65625 27285 65659 27319
rect 66269 27285 66303 27319
rect 66913 27285 66947 27319
rect 68201 27285 68235 27319
rect 68569 27285 68603 27319
rect 70041 27285 70075 27319
rect 70777 27285 70811 27319
rect 71145 27285 71179 27319
rect 71237 27285 71271 27319
rect 74273 27285 74307 27319
rect 75009 27285 75043 27319
rect 75101 27285 75135 27319
rect 75929 27285 75963 27319
rect 78689 27285 78723 27319
rect 79057 27285 79091 27319
rect 79885 27285 79919 27319
rect 83657 27285 83691 27319
rect 84485 27285 84519 27319
rect 88809 27285 88843 27319
rect 89821 27285 89855 27319
rect 90097 27285 90131 27319
rect 90465 27285 90499 27319
rect 91937 27285 91971 27319
rect 92857 27285 92891 27319
rect 94329 27285 94363 27319
rect 94697 27285 94731 27319
rect 95525 27285 95559 27319
rect 104817 27285 104851 27319
rect 105553 27285 105587 27319
rect 110061 27285 110095 27319
rect 112545 27285 112579 27319
rect 114569 27285 114603 27319
rect 116225 27285 116259 27319
rect 3341 27081 3375 27115
rect 4629 27081 4663 27115
rect 7849 27081 7883 27115
rect 10609 27081 10643 27115
rect 11713 27081 11747 27115
rect 27169 27081 27203 27115
rect 29377 27081 29411 27115
rect 32965 27081 32999 27115
rect 33885 27081 33919 27115
rect 35265 27081 35299 27115
rect 36461 27081 36495 27115
rect 38117 27081 38151 27115
rect 40509 27081 40543 27115
rect 41337 27081 41371 27115
rect 45845 27081 45879 27115
rect 52929 27081 52963 27115
rect 55321 27081 55355 27115
rect 56149 27081 56183 27115
rect 56517 27081 56551 27115
rect 57161 27081 57195 27115
rect 58357 27081 58391 27115
rect 58817 27081 58851 27115
rect 59185 27081 59219 27115
rect 77033 27081 77067 27115
rect 77401 27081 77435 27115
rect 79793 27081 79827 27115
rect 84761 27081 84795 27115
rect 90373 27081 90407 27115
rect 92857 27081 92891 27115
rect 94513 27081 94547 27115
rect 95709 27081 95743 27115
rect 100585 27081 100619 27115
rect 105369 27081 105403 27115
rect 111533 27081 111567 27115
rect 116317 27081 116351 27115
rect 15669 27013 15703 27047
rect 35633 27013 35667 27047
rect 46673 27013 46707 27047
rect 50721 27013 50755 27047
rect 53389 27013 53423 27047
rect 64889 27013 64923 27047
rect 68661 27013 68695 27047
rect 70317 27013 70351 27047
rect 76021 27013 76055 27047
rect 94421 27013 94455 27047
rect 104725 27013 104759 27047
rect 116777 27013 116811 27047
rect 117421 27013 117455 27047
rect 117697 27013 117731 27047
rect 1409 26945 1443 26979
rect 2881 26945 2915 26979
rect 3525 26945 3559 26979
rect 4813 26945 4847 26979
rect 8033 26945 8067 26979
rect 10793 26945 10827 26979
rect 11897 26945 11931 26979
rect 14289 26945 14323 26979
rect 14565 26945 14599 26979
rect 19901 26945 19935 26979
rect 20729 26945 20763 26979
rect 27353 26945 27387 26979
rect 29561 26945 29595 26979
rect 30389 26945 30423 26979
rect 33149 26945 33183 26979
rect 34069 26945 34103 26979
rect 34621 26945 34655 26979
rect 35725 26945 35759 26979
rect 36645 26945 36679 26979
rect 38301 26945 38335 26979
rect 40693 26945 40727 26979
rect 41521 26949 41555 26983
rect 46029 26945 46063 26979
rect 49525 26945 49559 26979
rect 50169 26945 50203 26979
rect 50905 26945 50939 26979
rect 51457 26945 51491 26979
rect 53113 26945 53147 26979
rect 55689 26945 55723 26979
rect 56333 26945 56367 26979
rect 56701 26945 56735 26979
rect 57345 26945 57379 26979
rect 59277 26945 59311 26979
rect 60013 26945 60047 26979
rect 61945 26945 61979 26979
rect 62589 26945 62623 26979
rect 63693 26945 63727 26979
rect 63785 26945 63819 26979
rect 65901 26945 65935 26979
rect 66545 26945 66579 26979
rect 69029 26945 69063 26979
rect 70133 26945 70167 26979
rect 70961 26945 70995 26979
rect 72249 26945 72283 26979
rect 73169 26945 73203 26979
rect 73629 26945 73663 26979
rect 74273 26945 74307 26979
rect 76665 26945 76699 26979
rect 77493 26945 77527 26979
rect 78137 26945 78171 26979
rect 78689 26945 78723 26979
rect 79333 26945 79367 26979
rect 79977 26945 80011 26979
rect 84081 26945 84115 26979
rect 84945 26945 84979 26979
rect 85589 26945 85623 26979
rect 86233 26945 86267 26979
rect 86877 26945 86911 26979
rect 89637 26945 89671 26979
rect 90281 26945 90315 26979
rect 91385 26945 91419 26979
rect 92397 26945 92431 26979
rect 93041 26945 93075 26979
rect 95249 26945 95283 26979
rect 95893 26945 95927 26979
rect 100769 26945 100803 26979
rect 103713 26945 103747 26979
rect 105553 26945 105587 26979
rect 111717 26945 111751 26979
rect 116501 26945 116535 26979
rect 117237 26945 117271 26979
rect 117973 26945 118007 26979
rect 1685 26877 1719 26911
rect 30481 26877 30515 26911
rect 30573 26877 30607 26911
rect 35909 26877 35943 26911
rect 39221 26877 39255 26911
rect 39497 26877 39531 26911
rect 48053 26877 48087 26911
rect 48329 26877 48363 26911
rect 51641 26877 51675 26911
rect 53665 26877 53699 26911
rect 53941 26877 53975 26911
rect 55781 26877 55815 26911
rect 55873 26877 55907 26911
rect 57897 26877 57931 26911
rect 59461 26877 59495 26911
rect 60289 26877 60323 26911
rect 62037 26877 62071 26911
rect 62221 26877 62255 26911
rect 63877 26877 63911 26911
rect 64981 26877 65015 26911
rect 65073 26877 65107 26911
rect 72341 26877 72375 26911
rect 72525 26877 72559 26911
rect 73353 26877 73387 26911
rect 76113 26877 76147 26911
rect 76205 26877 76239 26911
rect 77585 26877 77619 26911
rect 90557 26877 90591 26911
rect 2697 26809 2731 26843
rect 15853 26809 15887 26843
rect 20545 26809 20579 26843
rect 30021 26809 30055 26843
rect 49985 26809 50019 26843
rect 58173 26809 58207 26843
rect 65717 26809 65751 26843
rect 66361 26809 66395 26843
rect 71881 26809 71915 26843
rect 74503 26809 74537 26843
rect 79149 26809 79183 26843
rect 84301 26809 84335 26843
rect 86049 26809 86083 26843
rect 89913 26809 89947 26843
rect 92213 26809 92247 26843
rect 95065 26809 95099 26843
rect 104909 26809 104943 26843
rect 19993 26741 20027 26775
rect 34713 26741 34747 26775
rect 46949 26741 46983 26775
rect 49341 26741 49375 26775
rect 53481 26741 53515 26775
rect 61577 26741 61611 26775
rect 63325 26741 63359 26775
rect 64337 26741 64371 26775
rect 64521 26741 64555 26775
rect 70777 26741 70811 26775
rect 72985 26741 73019 26775
rect 75653 26741 75687 26775
rect 78505 26741 78539 26775
rect 85405 26741 85439 26775
rect 86693 26741 86727 26775
rect 89453 26741 89487 26775
rect 90925 26741 90959 26775
rect 91477 26741 91511 26775
rect 103529 26741 103563 26775
rect 118065 26741 118099 26775
rect 29745 26537 29779 26571
rect 46489 26537 46523 26571
rect 69121 26537 69155 26571
rect 70041 26537 70075 26571
rect 77401 26537 77435 26571
rect 2697 26469 2731 26503
rect 49065 26469 49099 26503
rect 53573 26469 53607 26503
rect 54585 26469 54619 26503
rect 55321 26469 55355 26503
rect 56425 26469 56459 26503
rect 58725 26469 58759 26503
rect 79149 26469 79183 26503
rect 117329 26469 117363 26503
rect 1409 26401 1443 26435
rect 35817 26401 35851 26435
rect 61853 26401 61887 26435
rect 79793 26401 79827 26435
rect 92029 26401 92063 26435
rect 1685 26333 1719 26367
rect 2881 26333 2915 26367
rect 29929 26333 29963 26367
rect 46673 26333 46707 26367
rect 48237 26333 48271 26367
rect 49249 26333 49283 26367
rect 50353 26333 50387 26367
rect 53757 26333 53791 26367
rect 54769 26333 54803 26367
rect 55505 26333 55539 26367
rect 56609 26333 56643 26367
rect 58909 26333 58943 26367
rect 62681 26333 62715 26367
rect 69305 26333 69339 26367
rect 70225 26333 70259 26367
rect 72065 26333 72099 26367
rect 75009 26333 75043 26367
rect 76481 26333 76515 26367
rect 77585 26333 77619 26367
rect 90465 26333 90499 26367
rect 93685 26333 93719 26367
rect 117145 26333 117179 26367
rect 117973 26333 118007 26367
rect 35633 26265 35667 26299
rect 61669 26265 61703 26299
rect 61761 26265 61795 26299
rect 71237 26265 71271 26299
rect 71421 26265 71455 26299
rect 79517 26265 79551 26299
rect 91845 26265 91879 26299
rect 118157 26265 118191 26299
rect 35173 26197 35207 26231
rect 35541 26197 35575 26231
rect 48053 26197 48087 26231
rect 50169 26197 50203 26231
rect 61301 26197 61335 26231
rect 62497 26197 62531 26231
rect 71881 26197 71915 26231
rect 74825 26197 74859 26231
rect 76665 26197 76699 26231
rect 79609 26197 79643 26231
rect 90281 26197 90315 26231
rect 93501 26197 93535 26231
rect 1409 25993 1443 26027
rect 35265 25993 35299 26027
rect 59921 25993 59955 26027
rect 61669 25993 61703 26027
rect 76113 25993 76147 26027
rect 117237 25993 117271 26027
rect 117973 25925 118007 25959
rect 1593 25857 1627 25891
rect 35449 25857 35483 25891
rect 57897 25857 57931 25891
rect 58081 25857 58115 25891
rect 60289 25857 60323 25891
rect 61853 25857 61887 25891
rect 76297 25857 76331 25891
rect 117421 25857 117455 25891
rect 60381 25789 60415 25823
rect 60565 25789 60599 25823
rect 118157 25721 118191 25755
rect 58265 25653 58299 25687
rect 58541 25653 58575 25687
rect 59553 25653 59587 25687
rect 32689 25381 32723 25415
rect 45109 25381 45143 25415
rect 58081 25381 58115 25415
rect 32873 25245 32907 25279
rect 45293 25245 45327 25279
rect 57897 25245 57931 25279
rect 64061 25245 64095 25279
rect 118157 25245 118191 25279
rect 36645 25177 36679 25211
rect 36829 25177 36863 25211
rect 64245 25177 64279 25211
rect 117973 25109 118007 25143
rect 31033 24905 31067 24939
rect 32137 24905 32171 24939
rect 1685 24769 1719 24803
rect 32505 24769 32539 24803
rect 118157 24769 118191 24803
rect 1409 24701 1443 24735
rect 31125 24701 31159 24735
rect 31309 24701 31343 24735
rect 32597 24701 32631 24735
rect 32781 24701 32815 24735
rect 33241 24701 33275 24735
rect 30665 24633 30699 24667
rect 31769 24565 31803 24599
rect 117605 24565 117639 24599
rect 117973 24565 118007 24599
rect 30665 24361 30699 24395
rect 31309 24225 31343 24259
rect 1409 24157 1443 24191
rect 1685 24157 1719 24191
rect 2881 24157 2915 24191
rect 30389 24089 30423 24123
rect 31033 24089 31067 24123
rect 2697 24021 2731 24055
rect 31125 24021 31159 24055
rect 1593 23681 1627 23715
rect 117605 23681 117639 23715
rect 117329 23613 117363 23647
rect 1409 23477 1443 23511
rect 94881 22661 94915 22695
rect 94789 22593 94823 22627
rect 95801 22593 95835 22627
rect 118157 22593 118191 22627
rect 94973 22525 95007 22559
rect 95433 22525 95467 22559
rect 94421 22457 94455 22491
rect 117973 22457 118007 22491
rect 95617 22389 95651 22423
rect 50721 22049 50755 22083
rect 1593 21981 1627 22015
rect 49525 21981 49559 22015
rect 50537 21981 50571 22015
rect 49341 21913 49375 21947
rect 68569 21913 68603 21947
rect 1409 21845 1443 21879
rect 50169 21845 50203 21879
rect 50629 21845 50663 21879
rect 68661 21845 68695 21879
rect 47777 21641 47811 21675
rect 68201 21641 68235 21675
rect 1409 21505 1443 21539
rect 47593 21505 47627 21539
rect 68569 21505 68603 21539
rect 68661 21437 68695 21471
rect 68753 21437 68787 21471
rect 117329 21437 117363 21471
rect 117605 21437 117639 21471
rect 1593 21301 1627 21335
rect 54677 21029 54711 21063
rect 72893 20961 72927 20995
rect 85037 20961 85071 20995
rect 54493 20893 54527 20927
rect 55781 20893 55815 20927
rect 72709 20893 72743 20927
rect 84853 20893 84887 20927
rect 118157 20893 118191 20927
rect 84209 20825 84243 20859
rect 84945 20825 84979 20859
rect 56057 20757 56091 20791
rect 72341 20757 72375 20791
rect 72801 20757 72835 20791
rect 84485 20757 84519 20791
rect 117973 20757 118007 20791
rect 79149 20553 79183 20587
rect 114569 20553 114603 20587
rect 71881 20417 71915 20451
rect 79057 20417 79091 20451
rect 79701 20417 79735 20451
rect 83657 20417 83691 20451
rect 114753 20417 114787 20451
rect 79241 20349 79275 20383
rect 83933 20349 83967 20383
rect 72065 20213 72099 20247
rect 78689 20213 78723 20247
rect 1593 19805 1627 19839
rect 80161 19805 80195 19839
rect 118157 19805 118191 19839
rect 79333 19737 79367 19771
rect 79517 19737 79551 19771
rect 113649 19737 113683 19771
rect 1409 19669 1443 19703
rect 79977 19669 80011 19703
rect 113741 19669 113775 19703
rect 117973 19669 118007 19703
rect 1869 19329 1903 19363
rect 2145 19125 2179 19159
rect 1593 18717 1627 18751
rect 117881 18717 117915 18751
rect 1409 18581 1443 18615
rect 118065 18581 118099 18615
rect 33333 18241 33367 18275
rect 117881 18241 117915 18275
rect 33057 18173 33091 18207
rect 118065 18037 118099 18071
rect 33333 17833 33367 17867
rect 33977 17697 34011 17731
rect 33701 17629 33735 17663
rect 33793 17493 33827 17527
rect 1593 17153 1627 17187
rect 82921 17153 82955 17187
rect 1409 17017 1443 17051
rect 1961 16949 1995 16983
rect 82737 16949 82771 16983
rect 81817 16677 81851 16711
rect 71513 16609 71547 16643
rect 82737 16609 82771 16643
rect 83289 16609 83323 16643
rect 117605 16609 117639 16643
rect 1593 16541 1627 16575
rect 66913 16541 66947 16575
rect 82645 16541 82679 16575
rect 117329 16541 117363 16575
rect 71237 16473 71271 16507
rect 82553 16473 82587 16507
rect 1409 16405 1443 16439
rect 67097 16405 67131 16439
rect 82185 16405 82219 16439
rect 68201 16133 68235 16167
rect 67005 16065 67039 16099
rect 68385 16065 68419 16099
rect 69305 16065 69339 16099
rect 66821 15929 66855 15963
rect 68569 15861 68603 15895
rect 69489 15861 69523 15895
rect 118157 15861 118191 15895
rect 69581 15657 69615 15691
rect 70777 15657 70811 15691
rect 66177 15521 66211 15555
rect 67281 15521 67315 15555
rect 67465 15521 67499 15555
rect 68293 15521 68327 15555
rect 71329 15521 71363 15555
rect 1593 15453 1627 15487
rect 64889 15453 64923 15487
rect 65993 15453 66027 15487
rect 67189 15453 67223 15487
rect 67373 15453 67407 15487
rect 68201 15453 68235 15487
rect 68385 15453 68419 15487
rect 68477 15453 68511 15487
rect 68937 15453 68971 15487
rect 69213 15453 69247 15487
rect 30665 15385 30699 15419
rect 30849 15385 30883 15419
rect 66085 15385 66119 15419
rect 66637 15385 66671 15419
rect 69397 15385 69431 15419
rect 1409 15317 1443 15351
rect 64705 15317 64739 15351
rect 65625 15317 65659 15351
rect 67005 15317 67039 15351
rect 68017 15317 68051 15351
rect 71145 15317 71179 15351
rect 71237 15317 71271 15351
rect 71881 15317 71915 15351
rect 10517 15113 10551 15147
rect 64245 15045 64279 15079
rect 65165 15045 65199 15079
rect 66545 15045 66579 15079
rect 67373 15045 67407 15079
rect 68753 15045 68787 15079
rect 69489 15045 69523 15079
rect 69765 15045 69799 15079
rect 8033 14977 8067 15011
rect 10701 14977 10735 15011
rect 49617 14977 49651 15011
rect 50445 14977 50479 15011
rect 53757 14977 53791 15011
rect 54861 14977 54895 15011
rect 55873 14977 55907 15011
rect 63969 14977 64003 15011
rect 64889 14977 64923 15011
rect 65901 14977 65935 15011
rect 67281 14977 67315 15011
rect 69213 14977 69247 15011
rect 69305 14977 69339 15011
rect 69949 14977 69983 15011
rect 70777 14977 70811 15011
rect 70961 14977 70995 15011
rect 50629 14909 50663 14943
rect 54585 14909 54619 14943
rect 56149 14909 56183 14943
rect 67557 14909 67591 14943
rect 70041 14909 70075 14943
rect 8217 14841 8251 14875
rect 66913 14841 66947 14875
rect 68753 14841 68787 14875
rect 49709 14773 49743 14807
rect 53849 14773 53883 14807
rect 65993 14773 66027 14807
rect 70133 14773 70167 14807
rect 70317 14773 70351 14807
rect 70869 14773 70903 14807
rect 55505 14569 55539 14603
rect 71605 14569 71639 14603
rect 118065 14569 118099 14603
rect 2237 14501 2271 14535
rect 66269 14433 66303 14467
rect 70849 14433 70883 14467
rect 1593 14365 1627 14399
rect 2421 14365 2455 14399
rect 50629 14365 50663 14399
rect 55321 14365 55355 14399
rect 64613 14365 64647 14399
rect 65993 14365 66027 14399
rect 66821 14365 66855 14399
rect 68661 14365 68695 14399
rect 71053 14365 71087 14399
rect 71513 14365 71547 14399
rect 117881 14365 117915 14399
rect 64889 14297 64923 14331
rect 67088 14297 67122 14331
rect 68928 14297 68962 14331
rect 70777 14297 70811 14331
rect 1409 14229 1443 14263
rect 50721 14229 50755 14263
rect 68201 14229 68235 14263
rect 70041 14229 70075 14263
rect 70961 14229 70995 14263
rect 65625 14025 65659 14059
rect 71237 14025 71271 14059
rect 85589 14025 85623 14059
rect 86233 14025 86267 14059
rect 118065 14025 118099 14059
rect 66536 13957 66570 13991
rect 65809 13889 65843 13923
rect 68569 13889 68603 13923
rect 107209 13889 107243 13923
rect 117881 13889 117915 13923
rect 66269 13821 66303 13855
rect 70777 13821 70811 13855
rect 86325 13821 86359 13855
rect 86417 13821 86451 13855
rect 107393 13821 107427 13855
rect 71053 13753 71087 13787
rect 67649 13685 67683 13719
rect 69857 13685 69891 13719
rect 85865 13685 85899 13719
rect 68937 13481 68971 13515
rect 70133 13481 70167 13515
rect 67649 13277 67683 13311
rect 70041 13277 70075 13311
rect 86785 13277 86819 13311
rect 118157 13277 118191 13311
rect 1869 13209 1903 13243
rect 1961 13141 1995 13175
rect 86601 13141 86635 13175
rect 117973 13141 118007 13175
rect 32137 12937 32171 12971
rect 67649 12937 67683 12971
rect 68201 12937 68235 12971
rect 69949 12937 69983 12971
rect 76757 12937 76791 12971
rect 66536 12869 66570 12903
rect 1593 12801 1627 12835
rect 32321 12801 32355 12835
rect 66269 12801 66303 12835
rect 68385 12801 68419 12835
rect 68477 12801 68511 12835
rect 69489 12801 69523 12835
rect 108221 12801 108255 12835
rect 68569 12733 68603 12767
rect 68661 12733 68695 12767
rect 76849 12733 76883 12767
rect 77033 12733 77067 12767
rect 76113 12665 76147 12699
rect 1409 12597 1443 12631
rect 69581 12597 69615 12631
rect 76389 12597 76423 12631
rect 108037 12597 108071 12631
rect 21465 12393 21499 12427
rect 31217 12393 31251 12427
rect 67281 12393 67315 12427
rect 67465 12393 67499 12427
rect 68293 12393 68327 12427
rect 22569 12257 22603 12291
rect 22753 12257 22787 12291
rect 31861 12257 31895 12291
rect 21649 12189 21683 12223
rect 31585 12189 31619 12223
rect 43729 12189 43763 12223
rect 67833 12189 67867 12223
rect 68201 12189 68235 12223
rect 22477 12121 22511 12155
rect 31677 12121 31711 12155
rect 44005 12121 44039 12155
rect 67097 12121 67131 12155
rect 67313 12121 67347 12155
rect 22109 12053 22143 12087
rect 30849 12053 30883 12087
rect 39221 11849 39255 11883
rect 76941 11781 76975 11815
rect 1593 11713 1627 11747
rect 39313 11645 39347 11679
rect 39405 11645 39439 11679
rect 117329 11645 117363 11679
rect 117605 11645 117639 11679
rect 1409 11577 1443 11611
rect 38485 11509 38519 11543
rect 38853 11509 38887 11543
rect 77033 11509 77067 11543
rect 117973 11237 118007 11271
rect 9229 11169 9263 11203
rect 42533 11169 42567 11203
rect 8953 11101 8987 11135
rect 42809 11101 42843 11135
rect 118157 11101 118191 11135
rect 66361 10761 66395 10795
rect 65073 10693 65107 10727
rect 1593 10625 1627 10659
rect 1409 10421 1443 10455
rect 2513 10217 2547 10251
rect 113741 10217 113775 10251
rect 2697 10013 2731 10047
rect 118157 10013 118191 10047
rect 1869 9945 1903 9979
rect 2053 9945 2087 9979
rect 113649 9945 113683 9979
rect 117973 9877 118007 9911
rect 114753 9537 114787 9571
rect 114569 9401 114603 9435
rect 1593 8449 1627 8483
rect 29745 8449 29779 8483
rect 117605 8449 117639 8483
rect 118157 8449 118191 8483
rect 29469 8381 29503 8415
rect 1409 8313 1443 8347
rect 117973 8313 118007 8347
rect 29745 8041 29779 8075
rect 77217 7973 77251 8007
rect 30297 7905 30331 7939
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 30113 7769 30147 7803
rect 77033 7769 77067 7803
rect 30205 7701 30239 7735
rect 30849 7701 30883 7735
rect 86233 7361 86267 7395
rect 117973 7361 118007 7395
rect 86325 7157 86359 7191
rect 118065 7157 118099 7191
rect 50353 6749 50387 6783
rect 50169 6613 50203 6647
rect 49893 6409 49927 6443
rect 1593 6273 1627 6307
rect 50261 6273 50295 6307
rect 50353 6273 50387 6307
rect 86969 6273 87003 6307
rect 117881 6273 117915 6307
rect 50445 6205 50479 6239
rect 1409 6137 1443 6171
rect 118065 6137 118099 6171
rect 1961 6069 1995 6103
rect 86785 6069 86819 6103
rect 1869 5593 1903 5627
rect 1961 5525 1995 5559
rect 83013 5253 83047 5287
rect 1409 5185 1443 5219
rect 82829 5185 82863 5219
rect 118157 5185 118191 5219
rect 1593 4981 1627 5015
rect 117973 4981 118007 5015
rect 79333 4573 79367 4607
rect 79793 4573 79827 4607
rect 79977 4505 80011 4539
rect 117789 4505 117823 4539
rect 117881 4437 117915 4471
rect 60657 4233 60691 4267
rect 82645 4233 82679 4267
rect 82553 4165 82587 4199
rect 117973 4165 118007 4199
rect 1593 4097 1627 4131
rect 59553 4097 59587 4131
rect 61025 4097 61059 4131
rect 62037 4097 62071 4131
rect 79241 4097 79275 4131
rect 116869 4097 116903 4131
rect 117421 4097 117455 4131
rect 60289 4029 60323 4063
rect 61117 4029 61151 4063
rect 61301 4029 61335 4063
rect 82737 4029 82771 4063
rect 1409 3961 1443 3995
rect 59369 3893 59403 3927
rect 61853 3893 61887 3927
rect 79057 3893 79091 3927
rect 82185 3893 82219 3927
rect 117237 3893 117271 3927
rect 118065 3893 118099 3927
rect 59645 3689 59679 3723
rect 40693 3621 40727 3655
rect 73997 3621 74031 3655
rect 118065 3621 118099 3655
rect 61117 3553 61151 3587
rect 1593 3485 1627 3519
rect 2237 3485 2271 3519
rect 2881 3485 2915 3519
rect 32873 3485 32907 3519
rect 40877 3485 40911 3519
rect 42809 3485 42843 3519
rect 46029 3485 46063 3519
rect 47041 3485 47075 3519
rect 47685 3485 47719 3519
rect 52469 3485 52503 3519
rect 57621 3485 57655 3519
rect 58257 3481 58291 3515
rect 70961 3485 70995 3519
rect 71605 3485 71639 3519
rect 72249 3485 72283 3519
rect 72617 3485 72651 3519
rect 73077 3485 73111 3519
rect 74181 3485 74215 3519
rect 75009 3485 75043 3519
rect 76113 3485 76147 3519
rect 116593 3485 116627 3519
rect 117421 3485 117455 3519
rect 117881 3485 117915 3519
rect 59553 3417 59587 3451
rect 60933 3417 60967 3451
rect 2053 3349 2087 3383
rect 2697 3349 2731 3383
rect 32689 3349 32723 3383
rect 42625 3349 42659 3383
rect 45845 3349 45879 3383
rect 46857 3349 46891 3383
rect 47501 3349 47535 3383
rect 57437 3349 57471 3383
rect 58081 3349 58115 3383
rect 70777 3349 70811 3383
rect 71421 3349 71455 3383
rect 72065 3349 72099 3383
rect 72893 3349 72927 3383
rect 74825 3349 74859 3383
rect 75929 3349 75963 3383
rect 116409 3349 116443 3383
rect 117237 3349 117271 3383
rect 2145 3145 2179 3179
rect 2513 3145 2547 3179
rect 10333 3145 10367 3179
rect 20729 3145 20763 3179
rect 28917 3145 28951 3179
rect 29653 3145 29687 3179
rect 41705 3145 41739 3179
rect 43085 3145 43119 3179
rect 43913 3145 43947 3179
rect 47777 3145 47811 3179
rect 58081 3145 58115 3179
rect 76941 3145 76975 3179
rect 117145 3145 117179 3179
rect 1869 3077 1903 3111
rect 32965 3077 32999 3111
rect 42993 3077 43027 3111
rect 45569 3077 45603 3111
rect 47041 3077 47075 3111
rect 56977 3077 57011 3111
rect 57069 3077 57103 3111
rect 60841 3077 60875 3111
rect 61025 3077 61059 3111
rect 70593 3077 70627 3111
rect 74549 3077 74583 3111
rect 75285 3077 75319 3111
rect 101321 3077 101355 3111
rect 107485 3077 107519 3111
rect 117053 3077 117087 3111
rect 2697 3009 2731 3043
rect 3065 3009 3099 3043
rect 3525 3009 3559 3043
rect 5457 3009 5491 3043
rect 6561 3009 6595 3043
rect 6929 3009 6963 3043
rect 7389 3009 7423 3043
rect 7849 3009 7883 3043
rect 10241 3009 10275 3043
rect 12265 3009 12299 3043
rect 14473 3009 14507 3043
rect 20913 3009 20947 3043
rect 24501 3009 24535 3043
rect 27629 3009 27663 3043
rect 28273 3009 28307 3043
rect 28733 3009 28767 3043
rect 29561 3009 29595 3043
rect 31585 3009 31619 3043
rect 32597 3009 32631 3043
rect 33609 3009 33643 3043
rect 35081 3009 35115 3043
rect 35541 3009 35575 3043
rect 36461 3009 36495 3043
rect 37657 3009 37691 3043
rect 38301 3009 38335 3043
rect 39589 3009 39623 3043
rect 40417 3009 40451 3043
rect 41889 3009 41923 3043
rect 44097 3009 44131 3043
rect 45385 3009 45419 3043
rect 46029 3009 46063 3043
rect 46857 3009 46891 3043
rect 47961 3009 47995 3043
rect 48605 3009 48639 3043
rect 51181 3009 51215 3043
rect 51917 3009 51951 3043
rect 53113 3009 53147 3043
rect 55689 3009 55723 3043
rect 57885 3009 57919 3043
rect 59001 3009 59035 3043
rect 59737 3009 59771 3043
rect 62129 3009 62163 3043
rect 64429 3009 64463 3043
rect 65257 3009 65291 3043
rect 66361 3009 66395 3043
rect 67005 3009 67039 3043
rect 68569 3009 68603 3043
rect 69857 3009 69891 3043
rect 70409 3009 70443 3043
rect 71237 3009 71271 3043
rect 72249 3009 72283 3043
rect 72341 3009 72375 3043
rect 73537 3009 73571 3043
rect 76849 3009 76883 3043
rect 77861 3009 77895 3043
rect 81449 3009 81483 3043
rect 87245 3009 87279 3043
rect 101505 3009 101539 3043
rect 102701 3009 102735 3043
rect 110337 3009 110371 3043
rect 111533 3009 111567 3043
rect 116225 3009 116259 3043
rect 117789 3009 117823 3043
rect 7573 2941 7607 2975
rect 37749 2941 37783 2975
rect 37841 2941 37875 2975
rect 40509 2941 40543 2975
rect 40693 2941 40727 2975
rect 43269 2941 43303 2975
rect 57253 2941 57287 2975
rect 59461 2941 59495 2975
rect 72433 2941 72467 2975
rect 77033 2941 77067 2975
rect 118065 2941 118099 2975
rect 3341 2873 3375 2907
rect 14289 2873 14323 2907
rect 27445 2873 27479 2907
rect 34897 2873 34931 2907
rect 35725 2873 35759 2907
rect 37289 2873 37323 2907
rect 52101 2873 52135 2907
rect 64613 2873 64647 2907
rect 66177 2873 66211 2907
rect 73353 2873 73387 2907
rect 76481 2873 76515 2907
rect 77677 2873 77711 2907
rect 107669 2873 107703 2907
rect 110153 2873 110187 2907
rect 111717 2873 111751 2907
rect 5273 2805 5307 2839
rect 6377 2805 6411 2839
rect 7205 2805 7239 2839
rect 12081 2805 12115 2839
rect 24317 2805 24351 2839
rect 26433 2805 26467 2839
rect 28089 2805 28123 2839
rect 31401 2805 31435 2839
rect 33425 2805 33459 2839
rect 36277 2805 36311 2839
rect 38117 2805 38151 2839
rect 39405 2805 39439 2839
rect 40049 2805 40083 2839
rect 42625 2805 42659 2839
rect 46213 2805 46247 2839
rect 48421 2805 48455 2839
rect 50997 2805 51031 2839
rect 52929 2805 52963 2839
rect 55505 2805 55539 2839
rect 56609 2805 56643 2839
rect 58817 2805 58851 2839
rect 61945 2805 61979 2839
rect 65073 2805 65107 2839
rect 66821 2805 66855 2839
rect 68385 2805 68419 2839
rect 69673 2805 69707 2839
rect 71329 2805 71363 2839
rect 71881 2805 71915 2839
rect 74641 2805 74675 2839
rect 75377 2805 75411 2839
rect 81265 2805 81299 2839
rect 87061 2805 87095 2839
rect 99297 2805 99331 2839
rect 102517 2805 102551 2839
rect 109785 2805 109819 2839
rect 116041 2805 116075 2839
rect 10885 2601 10919 2635
rect 14657 2601 14691 2635
rect 19809 2601 19843 2635
rect 22661 2601 22695 2635
rect 23305 2601 23339 2635
rect 25421 2601 25455 2635
rect 26985 2601 27019 2635
rect 28825 2601 28859 2635
rect 32137 2601 32171 2635
rect 58817 2601 58851 2635
rect 64521 2601 64555 2635
rect 66729 2601 66763 2635
rect 70777 2601 70811 2635
rect 71605 2601 71639 2635
rect 72617 2601 72651 2635
rect 82553 2601 82587 2635
rect 100217 2601 100251 2635
rect 100769 2601 100803 2635
rect 102241 2601 102275 2635
rect 103345 2601 103379 2635
rect 111073 2601 111107 2635
rect 114569 2601 114603 2635
rect 10241 2533 10275 2567
rect 11897 2533 11931 2567
rect 38485 2533 38519 2567
rect 47593 2533 47627 2567
rect 52745 2533 52779 2567
rect 54585 2533 54619 2567
rect 60657 2533 60691 2567
rect 68569 2533 68603 2567
rect 68937 2533 68971 2567
rect 69305 2533 69339 2567
rect 4905 2465 4939 2499
rect 27537 2465 27571 2499
rect 32781 2465 32815 2499
rect 34713 2465 34747 2499
rect 36645 2465 36679 2499
rect 40785 2465 40819 2499
rect 42441 2465 42475 2499
rect 46765 2465 46799 2499
rect 46949 2465 46983 2499
rect 48053 2465 48087 2499
rect 48237 2465 48271 2499
rect 52009 2465 52043 2499
rect 53205 2465 53239 2499
rect 53297 2465 53331 2499
rect 56793 2465 56827 2499
rect 59277 2465 59311 2499
rect 59461 2465 59495 2499
rect 61209 2465 61243 2499
rect 67281 2465 67315 2499
rect 69857 2465 69891 2499
rect 72065 2465 72099 2499
rect 72157 2465 72191 2499
rect 73997 2465 74031 2499
rect 77125 2465 77159 2499
rect 117881 2465 117915 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 2697 2397 2731 2431
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 9137 2397 9171 2431
rect 10425 2397 10459 2431
rect 11713 2397 11747 2431
rect 12633 2397 12667 2431
rect 15761 2397 15795 2431
rect 16865 2397 16899 2431
rect 17693 2397 17727 2431
rect 18337 2397 18371 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 20361 2397 20395 2431
rect 22201 2397 22235 2431
rect 22845 2397 22879 2431
rect 23489 2397 23523 2431
rect 24777 2397 24811 2431
rect 25237 2397 25271 2431
rect 26433 2397 26467 2431
rect 27353 2397 27387 2431
rect 27445 2397 27479 2431
rect 28365 2397 28399 2431
rect 29009 2397 29043 2431
rect 29929 2397 29963 2431
rect 30941 2397 30975 2431
rect 31585 2397 31619 2431
rect 33793 2397 33827 2431
rect 34989 2397 35023 2431
rect 36369 2397 36403 2431
rect 37657 2397 37691 2431
rect 38209 2397 38243 2431
rect 38669 2397 38703 2431
rect 39313 2397 39347 2431
rect 40509 2397 40543 2431
rect 42717 2397 42751 2431
rect 44465 2397 44499 2431
rect 46029 2397 46063 2431
rect 49249 2397 49283 2431
rect 50353 2397 50387 2431
rect 50997 2397 51031 2431
rect 54125 2397 54159 2431
rect 54769 2397 54803 2431
rect 56517 2397 56551 2431
rect 58173 2397 58207 2431
rect 62037 2397 62071 2431
rect 63417 2397 63451 2431
rect 64061 2397 64095 2431
rect 64705 2397 64739 2431
rect 65993 2397 66027 2431
rect 68017 2397 68051 2431
rect 69673 2397 69707 2431
rect 70961 2397 70995 2431
rect 73815 2397 73849 2431
rect 74457 2397 74491 2431
rect 75745 2397 75779 2431
rect 77953 2397 77987 2431
rect 78873 2397 78907 2431
rect 79517 2397 79551 2431
rect 81081 2397 81115 2431
rect 81357 2397 81391 2431
rect 82369 2397 82403 2431
rect 83657 2397 83691 2431
rect 84577 2397 84611 2431
rect 85313 2397 85347 2431
rect 86417 2397 86451 2431
rect 87429 2397 87463 2431
rect 87705 2397 87739 2431
rect 88993 2397 89027 2431
rect 89821 2397 89855 2431
rect 90465 2397 90499 2431
rect 91753 2397 91787 2431
rect 92397 2397 92431 2431
rect 92857 2397 92891 2431
rect 94329 2397 94363 2431
rect 95985 2397 96019 2431
rect 99757 2397 99791 2431
rect 100585 2397 100619 2431
rect 104633 2397 104667 2431
rect 106013 2397 106047 2431
rect 107025 2397 107059 2431
rect 107669 2397 107703 2431
rect 108313 2397 108347 2431
rect 110889 2397 110923 2431
rect 112177 2397 112211 2431
rect 112453 2397 112487 2431
rect 113649 2397 113683 2431
rect 114753 2397 114787 2431
rect 115397 2397 115431 2431
rect 3065 2329 3099 2363
rect 6745 2329 6779 2363
rect 10793 2329 10827 2363
rect 14565 2329 14599 2363
rect 32505 2329 32539 2363
rect 32597 2329 32631 2363
rect 33149 2329 33183 2363
rect 36461 2329 36495 2363
rect 41613 2329 41647 2363
rect 41797 2329 41831 2363
rect 45477 2329 45511 2363
rect 55873 2329 55907 2363
rect 59185 2329 59219 2363
rect 67097 2329 67131 2363
rect 76297 2329 76331 2363
rect 77033 2329 77067 2363
rect 94881 2329 94915 2363
rect 96997 2329 97031 2363
rect 98101 2329 98135 2363
rect 99573 2329 99607 2363
rect 102149 2329 102183 2363
rect 103253 2329 103287 2363
rect 105185 2329 105219 2363
rect 109877 2329 109911 2363
rect 116409 2329 116443 2363
rect 117605 2329 117639 2363
rect 7021 2261 7055 2295
rect 8217 2261 8251 2295
rect 8585 2261 8619 2295
rect 9321 2261 9355 2295
rect 9781 2261 9815 2295
rect 10149 2261 10183 2295
rect 12449 2261 12483 2295
rect 15577 2261 15611 2295
rect 16681 2261 16715 2295
rect 17509 2261 17543 2295
rect 18153 2261 18187 2295
rect 19257 2261 19291 2295
rect 24593 2261 24627 2295
rect 26249 2261 26283 2295
rect 28181 2261 28215 2295
rect 29745 2261 29779 2295
rect 30757 2261 30791 2295
rect 31401 2261 31435 2295
rect 33609 2261 33643 2295
rect 36001 2261 36035 2295
rect 37473 2261 37507 2295
rect 39129 2261 39163 2295
rect 40141 2261 40175 2295
rect 40601 2261 40635 2295
rect 41153 2261 41187 2295
rect 44281 2261 44315 2295
rect 45569 2261 45603 2295
rect 46305 2261 46339 2295
rect 46673 2261 46707 2295
rect 47961 2261 47995 2295
rect 49065 2261 49099 2295
rect 50169 2261 50203 2295
rect 50813 2261 50847 2295
rect 51457 2261 51491 2295
rect 51825 2261 51859 2295
rect 51917 2261 51951 2295
rect 53113 2261 53147 2295
rect 53941 2261 53975 2295
rect 55965 2261 55999 2295
rect 58265 2261 58299 2295
rect 61025 2261 61059 2295
rect 61117 2261 61151 2295
rect 61853 2261 61887 2295
rect 63233 2261 63267 2295
rect 63877 2261 63911 2295
rect 65809 2261 65843 2295
rect 66453 2261 66487 2295
rect 67189 2261 67223 2295
rect 67833 2261 67867 2295
rect 69765 2261 69799 2295
rect 70317 2261 70351 2295
rect 71237 2261 71271 2295
rect 71973 2261 72007 2295
rect 73629 2261 73663 2295
rect 74641 2261 74675 2295
rect 75561 2261 75595 2295
rect 76573 2261 76607 2295
rect 76941 2261 76975 2295
rect 77769 2261 77803 2295
rect 78689 2261 78723 2295
rect 79333 2261 79367 2295
rect 83841 2261 83875 2295
rect 84393 2261 84427 2295
rect 85129 2261 85163 2295
rect 86233 2261 86267 2295
rect 88809 2261 88843 2295
rect 89637 2261 89671 2295
rect 90281 2261 90315 2295
rect 91569 2261 91603 2295
rect 92213 2261 92247 2295
rect 93041 2261 93075 2295
rect 94145 2261 94179 2295
rect 94973 2261 95007 2295
rect 95801 2261 95835 2295
rect 97089 2261 97123 2295
rect 98193 2261 98227 2295
rect 104449 2261 104483 2295
rect 105277 2261 105311 2295
rect 105829 2261 105863 2295
rect 106841 2261 106875 2295
rect 107485 2261 107519 2295
rect 108129 2261 108163 2295
rect 109969 2261 110003 2295
rect 113465 2261 113499 2295
rect 115581 2261 115615 2295
rect 116501 2261 116535 2295
<< metal1 >>
rect 50798 28092 50804 28144
rect 50856 28132 50862 28144
rect 53098 28132 53104 28144
rect 50856 28104 53104 28132
rect 50856 28092 50862 28104
rect 53098 28092 53104 28104
rect 53156 28092 53162 28144
rect 40862 28024 40868 28076
rect 40920 28064 40926 28076
rect 46750 28064 46756 28076
rect 40920 28036 46756 28064
rect 40920 28024 40926 28036
rect 46750 28024 46756 28036
rect 46808 28024 46814 28076
rect 50706 28024 50712 28076
rect 50764 28064 50770 28076
rect 57606 28064 57612 28076
rect 50764 28036 57612 28064
rect 50764 28024 50770 28036
rect 57606 28024 57612 28036
rect 57664 28024 57670 28076
rect 69290 28024 69296 28076
rect 69348 28064 69354 28076
rect 75270 28064 75276 28076
rect 69348 28036 75276 28064
rect 69348 28024 69354 28036
rect 75270 28024 75276 28036
rect 75328 28024 75334 28076
rect 26694 27956 26700 28008
rect 26752 27996 26758 28008
rect 39574 27996 39580 28008
rect 26752 27968 39580 27996
rect 26752 27956 26758 27968
rect 39574 27956 39580 27968
rect 39632 27956 39638 28008
rect 39666 27956 39672 28008
rect 39724 27996 39730 28008
rect 40402 27996 40408 28008
rect 39724 27968 40408 27996
rect 39724 27956 39730 27968
rect 40402 27956 40408 27968
rect 40460 27996 40466 28008
rect 49142 27996 49148 28008
rect 40460 27968 49148 27996
rect 40460 27956 40466 27968
rect 49142 27956 49148 27968
rect 49200 27996 49206 28008
rect 49694 27996 49700 28008
rect 49200 27968 49700 27996
rect 49200 27956 49206 27968
rect 49694 27956 49700 27968
rect 49752 27956 49758 28008
rect 50246 27956 50252 28008
rect 50304 27996 50310 28008
rect 53466 27996 53472 28008
rect 50304 27968 53472 27996
rect 50304 27956 50310 27968
rect 53466 27956 53472 27968
rect 53524 27956 53530 28008
rect 59078 27956 59084 28008
rect 59136 27996 59142 28008
rect 62942 27996 62948 28008
rect 59136 27968 62948 27996
rect 59136 27956 59142 27968
rect 62942 27956 62948 27968
rect 63000 27956 63006 28008
rect 70302 27956 70308 28008
rect 70360 27996 70366 28008
rect 74994 27996 75000 28008
rect 70360 27968 75000 27996
rect 70360 27956 70366 27968
rect 74994 27956 75000 27968
rect 75052 27956 75058 28008
rect 40862 27928 40868 27940
rect 31864 27900 40868 27928
rect 9858 27820 9864 27872
rect 9916 27860 9922 27872
rect 17126 27860 17132 27872
rect 9916 27832 17132 27860
rect 9916 27820 9922 27832
rect 17126 27820 17132 27832
rect 17184 27820 17190 27872
rect 19794 27820 19800 27872
rect 19852 27860 19858 27872
rect 27062 27860 27068 27872
rect 19852 27832 27068 27860
rect 19852 27820 19858 27832
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 31754 27820 31760 27872
rect 31812 27860 31818 27872
rect 31864 27860 31892 27900
rect 40862 27888 40868 27900
rect 40920 27888 40926 27940
rect 40954 27888 40960 27940
rect 41012 27928 41018 27940
rect 41414 27928 41420 27940
rect 41012 27900 41420 27928
rect 41012 27888 41018 27900
rect 41414 27888 41420 27900
rect 41472 27888 41478 27940
rect 46474 27888 46480 27940
rect 46532 27928 46538 27940
rect 59722 27928 59728 27940
rect 46532 27900 59728 27928
rect 46532 27888 46538 27900
rect 59722 27888 59728 27900
rect 59780 27888 59786 27940
rect 61470 27888 61476 27940
rect 61528 27928 61534 27940
rect 68738 27928 68744 27940
rect 61528 27900 68744 27928
rect 61528 27888 61534 27900
rect 68738 27888 68744 27900
rect 68796 27928 68802 27940
rect 72878 27928 72884 27940
rect 68796 27900 72884 27928
rect 68796 27888 68802 27900
rect 72878 27888 72884 27900
rect 72936 27928 72942 27940
rect 76190 27928 76196 27940
rect 72936 27900 76196 27928
rect 72936 27888 72942 27900
rect 76190 27888 76196 27900
rect 76248 27888 76254 27940
rect 31812 27832 31892 27860
rect 31812 27820 31818 27832
rect 32674 27820 32680 27872
rect 32732 27860 32738 27872
rect 50798 27860 50804 27872
rect 32732 27832 50804 27860
rect 32732 27820 32738 27832
rect 50798 27820 50804 27832
rect 50856 27820 50862 27872
rect 50890 27820 50896 27872
rect 50948 27860 50954 27872
rect 54662 27860 54668 27872
rect 50948 27832 54668 27860
rect 50948 27820 50954 27832
rect 54662 27820 54668 27832
rect 54720 27820 54726 27872
rect 59354 27820 59360 27872
rect 59412 27860 59418 27872
rect 62114 27860 62120 27872
rect 59412 27832 62120 27860
rect 59412 27820 59418 27832
rect 62114 27820 62120 27832
rect 62172 27820 62178 27872
rect 68002 27820 68008 27872
rect 68060 27860 68066 27872
rect 68922 27860 68928 27872
rect 68060 27832 68928 27860
rect 68060 27820 68066 27832
rect 68922 27820 68928 27832
rect 68980 27820 68986 27872
rect 74442 27820 74448 27872
rect 74500 27860 74506 27872
rect 75914 27860 75920 27872
rect 74500 27832 75920 27860
rect 74500 27820 74506 27832
rect 75914 27820 75920 27832
rect 75972 27820 75978 27872
rect 78582 27820 78588 27872
rect 78640 27860 78646 27872
rect 79594 27860 79600 27872
rect 78640 27832 79600 27860
rect 78640 27820 78646 27832
rect 79594 27820 79600 27832
rect 79652 27820 79658 27872
rect 79778 27820 79784 27872
rect 79836 27860 79842 27872
rect 80422 27860 80428 27872
rect 79836 27832 80428 27860
rect 79836 27820 79842 27832
rect 80422 27820 80428 27832
rect 80480 27820 80486 27872
rect 84838 27820 84844 27872
rect 84896 27860 84902 27872
rect 93670 27860 93676 27872
rect 84896 27832 93676 27860
rect 84896 27820 84902 27832
rect 93670 27820 93676 27832
rect 93728 27820 93734 27872
rect 1104 27770 118864 27792
rect 1104 27718 15674 27770
rect 15726 27718 15738 27770
rect 15790 27718 15802 27770
rect 15854 27718 15866 27770
rect 15918 27718 15930 27770
rect 15982 27718 45122 27770
rect 45174 27718 45186 27770
rect 45238 27718 45250 27770
rect 45302 27718 45314 27770
rect 45366 27718 45378 27770
rect 45430 27718 74570 27770
rect 74622 27718 74634 27770
rect 74686 27718 74698 27770
rect 74750 27718 74762 27770
rect 74814 27718 74826 27770
rect 74878 27718 104018 27770
rect 104070 27718 104082 27770
rect 104134 27718 104146 27770
rect 104198 27718 104210 27770
rect 104262 27718 104274 27770
rect 104326 27718 118864 27770
rect 1104 27696 118864 27718
rect 17126 27616 17132 27668
rect 17184 27656 17190 27668
rect 84838 27656 84844 27668
rect 17184 27628 84844 27656
rect 17184 27616 17190 27628
rect 84838 27616 84844 27628
rect 84896 27616 84902 27668
rect 89714 27616 89720 27668
rect 89772 27656 89778 27668
rect 101674 27656 101680 27668
rect 89772 27628 95096 27656
rect 89772 27616 89778 27628
rect 9582 27588 9588 27600
rect 1596 27560 9588 27588
rect 1596 27461 1624 27560
rect 9582 27548 9588 27560
rect 9640 27548 9646 27600
rect 9677 27591 9735 27597
rect 9677 27557 9689 27591
rect 9723 27588 9735 27591
rect 9858 27588 9864 27600
rect 9723 27560 9864 27588
rect 9723 27557 9735 27560
rect 9677 27551 9735 27557
rect 9858 27548 9864 27560
rect 9916 27548 9922 27600
rect 10505 27591 10563 27597
rect 10505 27557 10517 27591
rect 10551 27588 10563 27591
rect 17034 27588 17040 27600
rect 10551 27560 17040 27588
rect 10551 27557 10563 27560
rect 10505 27551 10563 27557
rect 17034 27548 17040 27560
rect 17092 27548 17098 27600
rect 18690 27548 18696 27600
rect 18748 27588 18754 27600
rect 19245 27591 19303 27597
rect 19245 27588 19257 27591
rect 18748 27560 19257 27588
rect 18748 27548 18754 27560
rect 19245 27557 19257 27560
rect 19291 27557 19303 27591
rect 19245 27551 19303 27557
rect 19334 27548 19340 27600
rect 19392 27588 19398 27600
rect 22646 27588 22652 27600
rect 19392 27560 22508 27588
rect 22607 27560 22652 27588
rect 19392 27548 19398 27560
rect 2406 27520 2412 27532
rect 2367 27492 2412 27520
rect 2406 27480 2412 27492
rect 2464 27480 2470 27532
rect 4982 27520 4988 27532
rect 4943 27492 4988 27520
rect 4982 27480 4988 27492
rect 5040 27480 5046 27532
rect 6362 27520 6368 27532
rect 6323 27492 6368 27520
rect 6362 27480 6368 27492
rect 6420 27480 6426 27532
rect 7561 27523 7619 27529
rect 7561 27489 7573 27523
rect 7607 27520 7619 27523
rect 8113 27523 8171 27529
rect 8113 27520 8125 27523
rect 7607 27492 8125 27520
rect 7607 27489 7619 27492
rect 7561 27483 7619 27489
rect 8113 27489 8125 27492
rect 8159 27520 8171 27523
rect 22370 27520 22376 27532
rect 8159 27492 22376 27520
rect 8159 27489 8171 27492
rect 8113 27483 8171 27489
rect 22370 27480 22376 27492
rect 22428 27480 22434 27532
rect 22480 27520 22508 27560
rect 22646 27548 22652 27560
rect 22704 27548 22710 27600
rect 27154 27588 27160 27600
rect 23492 27560 27160 27588
rect 23382 27520 23388 27532
rect 22480 27492 23388 27520
rect 23382 27480 23388 27492
rect 23440 27480 23446 27532
rect 1581 27455 1639 27461
rect 1581 27421 1593 27455
rect 1627 27421 1639 27455
rect 2682 27452 2688 27464
rect 2643 27424 2688 27452
rect 1581 27415 1639 27421
rect 2682 27412 2688 27424
rect 2740 27412 2746 27464
rect 3602 27412 3608 27464
rect 3660 27452 3666 27464
rect 4249 27455 4307 27461
rect 4249 27452 4261 27455
rect 3660 27424 4261 27452
rect 3660 27412 3666 27424
rect 4249 27421 4261 27424
rect 4295 27421 4307 27455
rect 4249 27415 4307 27421
rect 5261 27455 5319 27461
rect 5261 27421 5273 27455
rect 5307 27421 5319 27455
rect 6638 27452 6644 27464
rect 6599 27424 6644 27452
rect 5261 27415 5319 27421
rect 4430 27384 4436 27396
rect 4391 27356 4436 27384
rect 4430 27344 4436 27356
rect 4488 27344 4494 27396
rect 1394 27316 1400 27328
rect 1355 27288 1400 27316
rect 1394 27276 1400 27288
rect 1452 27276 1458 27328
rect 5276 27316 5304 27415
rect 6638 27412 6644 27424
rect 6696 27412 6702 27464
rect 7098 27412 7104 27464
rect 7156 27452 7162 27464
rect 7929 27455 7987 27461
rect 7929 27452 7941 27455
rect 7156 27424 7941 27452
rect 7156 27412 7162 27424
rect 7929 27421 7941 27424
rect 7975 27421 7987 27455
rect 7929 27415 7987 27421
rect 11054 27412 11060 27464
rect 11112 27452 11118 27464
rect 11609 27455 11667 27461
rect 11609 27452 11621 27455
rect 11112 27424 11621 27452
rect 11112 27412 11118 27424
rect 11609 27421 11621 27424
rect 11655 27421 11667 27455
rect 11609 27415 11667 27421
rect 12434 27412 12440 27464
rect 12492 27452 12498 27464
rect 12492 27424 12537 27452
rect 12492 27412 12498 27424
rect 13814 27412 13820 27464
rect 13872 27452 13878 27464
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 13872 27424 14289 27452
rect 13872 27412 13878 27424
rect 14277 27421 14289 27424
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 15289 27455 15347 27461
rect 15289 27421 15301 27455
rect 15335 27421 15347 27455
rect 15289 27415 15347 27421
rect 15565 27455 15623 27461
rect 15565 27421 15577 27455
rect 15611 27452 15623 27455
rect 16022 27452 16028 27464
rect 15611 27424 16028 27452
rect 15611 27421 15623 27424
rect 15565 27415 15623 27421
rect 9398 27384 9404 27396
rect 9359 27356 9404 27384
rect 9398 27344 9404 27356
rect 9456 27344 9462 27396
rect 10318 27384 10324 27396
rect 10279 27356 10324 27384
rect 10318 27344 10324 27356
rect 10376 27344 10382 27396
rect 11149 27387 11207 27393
rect 11149 27353 11161 27387
rect 11195 27384 11207 27387
rect 11793 27387 11851 27393
rect 11793 27384 11805 27387
rect 11195 27356 11805 27384
rect 11195 27353 11207 27356
rect 11149 27347 11207 27353
rect 11793 27353 11805 27356
rect 11839 27384 11851 27387
rect 12161 27387 12219 27393
rect 12161 27384 12173 27387
rect 11839 27356 12173 27384
rect 11839 27353 11851 27356
rect 11793 27347 11851 27353
rect 12161 27353 12173 27356
rect 12207 27384 12219 27387
rect 15194 27384 15200 27396
rect 12207 27356 15200 27384
rect 12207 27353 12219 27356
rect 12161 27347 12219 27353
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 15304 27384 15332 27415
rect 16022 27412 16028 27424
rect 16080 27412 16086 27464
rect 17218 27452 17224 27464
rect 17179 27424 17224 27452
rect 17218 27412 17224 27424
rect 17276 27412 17282 27464
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27452 17923 27455
rect 18046 27452 18052 27464
rect 17911 27424 18052 27452
rect 17911 27421 17923 27424
rect 17865 27415 17923 27421
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27421 19487 27455
rect 20162 27452 20168 27464
rect 20123 27424 20168 27452
rect 19429 27415 19487 27421
rect 16114 27384 16120 27396
rect 15304 27356 16120 27384
rect 16114 27344 16120 27356
rect 16172 27344 16178 27396
rect 16206 27344 16212 27396
rect 16264 27384 16270 27396
rect 19334 27384 19340 27396
rect 16264 27356 19340 27384
rect 16264 27344 16270 27356
rect 19334 27344 19340 27356
rect 19392 27344 19398 27396
rect 19444 27384 19472 27415
rect 20162 27412 20168 27424
rect 20220 27412 20226 27464
rect 20346 27452 20352 27464
rect 20307 27424 20352 27452
rect 20346 27412 20352 27424
rect 20404 27412 20410 27464
rect 20530 27412 20536 27464
rect 20588 27452 20594 27464
rect 20993 27455 21051 27461
rect 20993 27452 21005 27455
rect 20588 27424 21005 27452
rect 20588 27412 20594 27424
rect 20993 27421 21005 27424
rect 21039 27421 21051 27455
rect 20993 27415 21051 27421
rect 21082 27412 21088 27464
rect 21140 27452 21146 27464
rect 21140 27424 22048 27452
rect 21140 27412 21146 27424
rect 21910 27384 21916 27396
rect 19444 27356 21916 27384
rect 21910 27344 21916 27356
rect 21968 27344 21974 27396
rect 22020 27384 22048 27424
rect 22094 27412 22100 27464
rect 22152 27452 22158 27464
rect 22189 27455 22247 27461
rect 22189 27452 22201 27455
rect 22152 27424 22201 27452
rect 22152 27412 22158 27424
rect 22189 27421 22201 27424
rect 22235 27421 22247 27455
rect 22189 27415 22247 27421
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 23492 27452 23520 27560
rect 27154 27548 27160 27560
rect 27212 27548 27218 27600
rect 31386 27588 31392 27600
rect 27356 27560 31392 27588
rect 23566 27480 23572 27532
rect 23624 27520 23630 27532
rect 23624 27492 27108 27520
rect 23624 27480 23630 27492
rect 23658 27452 23664 27464
rect 22879 27424 23520 27452
rect 23584 27424 23664 27452
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 23584 27384 23612 27424
rect 23658 27412 23664 27424
rect 23716 27412 23722 27464
rect 23842 27452 23848 27464
rect 23803 27424 23848 27452
rect 23842 27412 23848 27424
rect 23900 27412 23906 27464
rect 24581 27455 24639 27461
rect 24581 27421 24593 27455
rect 24627 27452 24639 27455
rect 25130 27452 25136 27464
rect 24627 27424 25136 27452
rect 24627 27421 24639 27424
rect 24581 27415 24639 27421
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 25314 27452 25320 27464
rect 25275 27424 25320 27452
rect 25314 27412 25320 27424
rect 25372 27412 25378 27464
rect 26418 27412 26424 27464
rect 26476 27452 26482 27464
rect 26973 27455 27031 27461
rect 26973 27452 26985 27455
rect 26476 27424 26985 27452
rect 26476 27412 26482 27424
rect 26973 27421 26985 27424
rect 27019 27421 27031 27455
rect 27080 27452 27108 27492
rect 27356 27452 27384 27560
rect 31386 27548 31392 27560
rect 31444 27548 31450 27600
rect 31754 27588 31760 27600
rect 31496 27560 31760 27588
rect 30650 27520 30656 27532
rect 27080 27424 27384 27452
rect 27724 27492 30656 27520
rect 26973 27415 27031 27421
rect 26878 27384 26884 27396
rect 22020 27356 23612 27384
rect 24320 27356 26884 27384
rect 11974 27316 11980 27328
rect 5276 27288 11980 27316
rect 11974 27276 11980 27288
rect 12032 27276 12038 27328
rect 12526 27316 12532 27328
rect 12487 27288 12532 27316
rect 12526 27276 12532 27288
rect 12584 27276 12590 27328
rect 14093 27319 14151 27325
rect 14093 27285 14105 27319
rect 14139 27316 14151 27319
rect 17126 27316 17132 27328
rect 14139 27288 17132 27316
rect 14139 27285 14151 27288
rect 14093 27279 14151 27285
rect 17126 27276 17132 27288
rect 17184 27276 17190 27328
rect 17310 27316 17316 27328
rect 17271 27288 17316 27316
rect 17310 27276 17316 27288
rect 17368 27276 17374 27328
rect 18095 27319 18153 27325
rect 18095 27285 18107 27319
rect 18141 27316 18153 27319
rect 20622 27316 20628 27328
rect 18141 27288 20628 27316
rect 18141 27285 18153 27288
rect 18095 27279 18153 27285
rect 20622 27276 20628 27288
rect 20680 27276 20686 27328
rect 20806 27316 20812 27328
rect 20767 27288 20812 27316
rect 20806 27276 20812 27288
rect 20864 27276 20870 27328
rect 22002 27316 22008 27328
rect 21963 27288 22008 27316
rect 22002 27276 22008 27288
rect 22060 27276 22066 27328
rect 22278 27276 22284 27328
rect 22336 27316 22342 27328
rect 23566 27316 23572 27328
rect 22336 27288 23572 27316
rect 22336 27276 22342 27288
rect 23566 27276 23572 27288
rect 23624 27276 23630 27328
rect 23661 27319 23719 27325
rect 23661 27285 23673 27319
rect 23707 27316 23719 27319
rect 24320 27316 24348 27356
rect 26878 27344 26884 27356
rect 26936 27344 26942 27396
rect 27522 27384 27528 27396
rect 26988 27356 27528 27384
rect 26988 27328 27016 27356
rect 27522 27344 27528 27356
rect 27580 27344 27586 27396
rect 23707 27288 24348 27316
rect 23707 27285 23719 27288
rect 23661 27279 23719 27285
rect 24394 27276 24400 27328
rect 24452 27316 24458 27328
rect 24949 27319 25007 27325
rect 24452 27288 24497 27316
rect 24452 27276 24458 27288
rect 24949 27285 24961 27319
rect 24995 27316 25007 27319
rect 25409 27319 25467 27325
rect 25409 27316 25421 27319
rect 24995 27288 25421 27316
rect 24995 27285 25007 27288
rect 24949 27279 25007 27285
rect 25409 27285 25421 27288
rect 25455 27316 25467 27319
rect 25869 27319 25927 27325
rect 25869 27316 25881 27319
rect 25455 27288 25881 27316
rect 25455 27285 25467 27288
rect 25409 27279 25467 27285
rect 25869 27285 25881 27288
rect 25915 27316 25927 27319
rect 26694 27316 26700 27328
rect 25915 27288 26700 27316
rect 25915 27285 25927 27288
rect 25869 27279 25927 27285
rect 26694 27276 26700 27288
rect 26752 27276 26758 27328
rect 26970 27276 26976 27328
rect 27028 27276 27034 27328
rect 27157 27319 27215 27325
rect 27157 27285 27169 27319
rect 27203 27316 27215 27319
rect 27724 27316 27752 27492
rect 30650 27480 30656 27492
rect 30708 27480 30714 27532
rect 30742 27480 30748 27532
rect 30800 27520 30806 27532
rect 30800 27492 30845 27520
rect 30800 27480 30806 27492
rect 31110 27480 31116 27532
rect 31168 27520 31174 27532
rect 31496 27520 31524 27560
rect 31754 27548 31760 27560
rect 31812 27548 31818 27600
rect 33042 27588 33048 27600
rect 31956 27560 33048 27588
rect 31846 27520 31852 27532
rect 31168 27492 31524 27520
rect 31726 27492 31852 27520
rect 31168 27480 31174 27492
rect 28074 27452 28080 27464
rect 28035 27424 28080 27452
rect 28074 27412 28080 27424
rect 28132 27412 28138 27464
rect 28813 27455 28871 27461
rect 28813 27421 28825 27455
rect 28859 27452 28871 27455
rect 28902 27452 28908 27464
rect 28859 27424 28908 27452
rect 28859 27421 28871 27424
rect 28813 27415 28871 27421
rect 28902 27412 28908 27424
rect 28960 27412 28966 27464
rect 30469 27455 30527 27461
rect 29380 27424 30420 27452
rect 29380 27384 29408 27424
rect 30282 27384 30288 27396
rect 27908 27356 29408 27384
rect 29472 27356 30288 27384
rect 27908 27325 27936 27356
rect 27203 27288 27752 27316
rect 27893 27319 27951 27325
rect 27203 27285 27215 27288
rect 27157 27279 27215 27285
rect 27893 27285 27905 27319
rect 27939 27285 27951 27319
rect 27893 27279 27951 27285
rect 28445 27319 28503 27325
rect 28445 27285 28457 27319
rect 28491 27316 28503 27319
rect 28905 27319 28963 27325
rect 28905 27316 28917 27319
rect 28491 27288 28917 27316
rect 28491 27285 28503 27288
rect 28445 27279 28503 27285
rect 28905 27285 28917 27288
rect 28951 27316 28963 27319
rect 29472 27316 29500 27356
rect 30282 27344 30288 27356
rect 30340 27344 30346 27396
rect 30392 27384 30420 27424
rect 30469 27421 30481 27455
rect 30515 27452 30527 27455
rect 30834 27452 30840 27464
rect 30515 27424 30840 27452
rect 30515 27421 30527 27424
rect 30469 27415 30527 27421
rect 30834 27412 30840 27424
rect 30892 27412 30898 27464
rect 30926 27412 30932 27464
rect 30984 27452 30990 27464
rect 31389 27455 31447 27461
rect 31389 27452 31401 27455
rect 30984 27424 31401 27452
rect 30984 27412 30990 27424
rect 31389 27421 31401 27424
rect 31435 27421 31447 27455
rect 31726 27452 31754 27492
rect 31846 27480 31852 27492
rect 31904 27480 31910 27532
rect 31389 27415 31447 27421
rect 31496 27424 31754 27452
rect 31956 27448 31984 27560
rect 33042 27548 33048 27560
rect 33100 27548 33106 27600
rect 33152 27560 34836 27588
rect 32030 27480 32036 27532
rect 32088 27520 32094 27532
rect 33152 27520 33180 27560
rect 33318 27520 33324 27532
rect 32088 27492 33180 27520
rect 33279 27492 33324 27520
rect 32088 27480 32094 27492
rect 33318 27480 33324 27492
rect 33376 27480 33382 27532
rect 34698 27520 34704 27532
rect 33428 27492 33732 27520
rect 34659 27492 34704 27520
rect 32585 27455 32643 27461
rect 32585 27452 32597 27455
rect 31496 27384 31524 27424
rect 31864 27420 31984 27448
rect 32048 27424 32597 27452
rect 30392 27356 31524 27384
rect 31570 27344 31576 27396
rect 31628 27384 31634 27396
rect 31864 27384 31892 27420
rect 32048 27396 32076 27424
rect 32585 27421 32597 27424
rect 32631 27421 32643 27455
rect 33428 27452 33456 27492
rect 33594 27452 33600 27464
rect 32585 27415 32643 27421
rect 32692 27424 33456 27452
rect 33555 27424 33600 27452
rect 31628 27356 31892 27384
rect 31628 27344 31634 27356
rect 32030 27344 32036 27396
rect 32088 27344 32094 27396
rect 32122 27344 32128 27396
rect 32180 27384 32186 27396
rect 32692 27384 32720 27424
rect 33594 27412 33600 27424
rect 33652 27412 33658 27464
rect 33704 27452 33732 27492
rect 34698 27480 34704 27492
rect 34756 27480 34762 27532
rect 34808 27520 34836 27560
rect 34882 27548 34888 27600
rect 34940 27588 34946 27600
rect 38194 27588 38200 27600
rect 34940 27560 38200 27588
rect 34940 27548 34946 27560
rect 38194 27548 38200 27560
rect 38252 27548 38258 27600
rect 39117 27591 39175 27597
rect 39117 27557 39129 27591
rect 39163 27588 39175 27591
rect 39942 27588 39948 27600
rect 39163 27560 39948 27588
rect 39163 27557 39175 27560
rect 39117 27551 39175 27557
rect 39942 27548 39948 27560
rect 40000 27548 40006 27600
rect 40586 27588 40592 27600
rect 40236 27560 40592 27588
rect 40236 27520 40264 27560
rect 40586 27548 40592 27560
rect 40644 27548 40650 27600
rect 40678 27548 40684 27600
rect 40736 27588 40742 27600
rect 40736 27560 42748 27588
rect 40736 27548 40742 27560
rect 40402 27520 40408 27532
rect 34808 27492 40264 27520
rect 40363 27492 40408 27520
rect 40402 27480 40408 27492
rect 40460 27480 40466 27532
rect 41230 27480 41236 27532
rect 41288 27520 41294 27532
rect 41693 27523 41751 27529
rect 41693 27520 41705 27523
rect 41288 27492 41705 27520
rect 41288 27480 41294 27492
rect 41693 27489 41705 27492
rect 41739 27489 41751 27523
rect 42720 27520 42748 27560
rect 42794 27548 42800 27600
rect 42852 27588 42858 27600
rect 43165 27591 43223 27597
rect 43165 27588 43177 27591
rect 42852 27560 43177 27588
rect 42852 27548 42858 27560
rect 43165 27557 43177 27560
rect 43211 27557 43223 27591
rect 43165 27551 43223 27557
rect 43901 27591 43959 27597
rect 43901 27557 43913 27591
rect 43947 27557 43959 27591
rect 43901 27551 43959 27557
rect 45005 27591 45063 27597
rect 45005 27557 45017 27591
rect 45051 27588 45063 27591
rect 50522 27588 50528 27600
rect 45051 27560 50528 27588
rect 45051 27557 45063 27560
rect 45005 27551 45063 27557
rect 43806 27520 43812 27532
rect 42720 27492 43812 27520
rect 41693 27483 41751 27489
rect 43806 27480 43812 27492
rect 43864 27480 43870 27532
rect 43916 27520 43944 27551
rect 50522 27548 50528 27560
rect 50580 27548 50586 27600
rect 53466 27588 53472 27600
rect 53427 27560 53472 27588
rect 53466 27548 53472 27560
rect 53524 27548 53530 27600
rect 54110 27548 54116 27600
rect 54168 27588 54174 27600
rect 59354 27588 59360 27600
rect 54168 27560 59360 27588
rect 54168 27548 54174 27560
rect 59354 27548 59360 27560
rect 59412 27548 59418 27600
rect 59446 27548 59452 27600
rect 59504 27588 59510 27600
rect 61102 27588 61108 27600
rect 59504 27560 61108 27588
rect 59504 27548 59510 27560
rect 61102 27548 61108 27560
rect 61160 27548 61166 27600
rect 61194 27548 61200 27600
rect 61252 27588 61258 27600
rect 61841 27591 61899 27597
rect 61841 27588 61853 27591
rect 61252 27560 61853 27588
rect 61252 27548 61258 27560
rect 61841 27557 61853 27560
rect 61887 27557 61899 27591
rect 61841 27551 61899 27557
rect 61948 27560 68968 27588
rect 43916 27492 49096 27520
rect 34882 27452 34888 27464
rect 33704 27424 34888 27452
rect 34882 27412 34888 27424
rect 34940 27412 34946 27464
rect 34977 27455 35035 27461
rect 34977 27421 34989 27455
rect 35023 27452 35035 27455
rect 35066 27452 35072 27464
rect 35023 27424 35072 27452
rect 35023 27421 35035 27424
rect 34977 27415 35035 27421
rect 35066 27412 35072 27424
rect 35124 27412 35130 27464
rect 35897 27455 35955 27461
rect 35897 27421 35909 27455
rect 35943 27452 35955 27455
rect 36449 27455 36507 27461
rect 36449 27452 36461 27455
rect 35943 27424 36461 27452
rect 35943 27421 35955 27424
rect 35897 27415 35955 27421
rect 36449 27421 36461 27424
rect 36495 27452 36507 27455
rect 36495 27424 36768 27452
rect 36495 27421 36507 27424
rect 36449 27415 36507 27421
rect 32180 27356 32720 27384
rect 32180 27344 32186 27356
rect 32766 27344 32772 27396
rect 32824 27384 32830 27396
rect 32824 27356 32869 27384
rect 32824 27344 32830 27356
rect 36262 27344 36268 27396
rect 36320 27384 36326 27396
rect 36740 27393 36768 27424
rect 37366 27412 37372 27464
rect 37424 27452 37430 27464
rect 37737 27455 37795 27461
rect 37737 27452 37749 27455
rect 37424 27424 37749 27452
rect 37424 27412 37430 27424
rect 37737 27421 37749 27424
rect 37783 27421 37795 27455
rect 37737 27415 37795 27421
rect 38657 27455 38715 27461
rect 38657 27421 38669 27455
rect 38703 27452 38715 27455
rect 39206 27452 39212 27464
rect 38703 27424 39212 27452
rect 38703 27421 38715 27424
rect 38657 27415 38715 27421
rect 39206 27412 39212 27424
rect 39264 27412 39270 27464
rect 39301 27455 39359 27461
rect 39301 27421 39313 27455
rect 39347 27452 39359 27455
rect 40494 27452 40500 27464
rect 39347 27424 40500 27452
rect 39347 27421 39359 27424
rect 39301 27415 39359 27421
rect 40494 27412 40500 27424
rect 40552 27412 40558 27464
rect 40586 27412 40592 27464
rect 40644 27452 40650 27464
rect 41509 27455 41567 27461
rect 41509 27452 41521 27455
rect 40644 27424 41521 27452
rect 40644 27412 40650 27424
rect 41509 27421 41521 27424
rect 41555 27421 41567 27455
rect 41509 27415 41567 27421
rect 41874 27412 41880 27464
rect 41932 27452 41938 27464
rect 42429 27455 42487 27461
rect 42429 27452 42441 27455
rect 41932 27424 42441 27452
rect 41932 27412 41938 27424
rect 42429 27421 42441 27424
rect 42475 27421 42487 27455
rect 43346 27452 43352 27464
rect 43307 27424 43352 27452
rect 42429 27415 42487 27421
rect 43346 27412 43352 27424
rect 43404 27412 43410 27464
rect 44082 27452 44088 27464
rect 44043 27424 44088 27452
rect 44082 27412 44088 27424
rect 44140 27412 44146 27464
rect 44450 27412 44456 27464
rect 44508 27452 44514 27464
rect 45189 27455 45247 27461
rect 45189 27452 45201 27455
rect 44508 27424 45201 27452
rect 44508 27412 44514 27424
rect 45189 27421 45201 27424
rect 45235 27421 45247 27455
rect 45189 27415 45247 27421
rect 47029 27455 47087 27461
rect 47029 27421 47041 27455
rect 47075 27452 47087 27455
rect 47210 27452 47216 27464
rect 47075 27424 47216 27452
rect 47075 27421 47087 27424
rect 47029 27415 47087 27421
rect 47210 27412 47216 27424
rect 47268 27412 47274 27464
rect 48133 27455 48191 27461
rect 48133 27421 48145 27455
rect 48179 27452 48191 27455
rect 48314 27452 48320 27464
rect 48179 27424 48320 27452
rect 48179 27421 48191 27424
rect 48133 27415 48191 27421
rect 48314 27412 48320 27424
rect 48372 27412 48378 27464
rect 49068 27452 49096 27492
rect 49142 27480 49148 27532
rect 49200 27520 49206 27532
rect 49329 27523 49387 27529
rect 49329 27520 49341 27523
rect 49200 27492 49341 27520
rect 49200 27480 49206 27492
rect 49329 27489 49341 27492
rect 49375 27489 49387 27523
rect 53484 27520 53512 27548
rect 54297 27523 54355 27529
rect 54297 27520 54309 27523
rect 53484 27492 54309 27520
rect 49329 27483 49387 27489
rect 54297 27489 54309 27492
rect 54343 27489 54355 27523
rect 54297 27483 54355 27489
rect 54478 27480 54484 27532
rect 54536 27520 54542 27532
rect 54536 27492 54581 27520
rect 54536 27480 54542 27492
rect 54662 27480 54668 27532
rect 54720 27520 54726 27532
rect 60734 27520 60740 27532
rect 54720 27492 60740 27520
rect 54720 27480 54726 27492
rect 60734 27480 60740 27492
rect 60792 27480 60798 27532
rect 60918 27480 60924 27532
rect 60976 27520 60982 27532
rect 61948 27520 61976 27560
rect 62114 27520 62120 27532
rect 60976 27492 61976 27520
rect 62040 27492 62120 27520
rect 60976 27480 60982 27492
rect 49068 27424 49280 27452
rect 36725 27387 36783 27393
rect 36320 27356 36365 27384
rect 36320 27344 36326 27356
rect 36725 27353 36737 27387
rect 36771 27384 36783 27387
rect 37642 27384 37648 27396
rect 36771 27356 37648 27384
rect 36771 27353 36783 27356
rect 36725 27347 36783 27353
rect 37642 27344 37648 27356
rect 37700 27344 37706 27396
rect 37918 27344 37924 27396
rect 37976 27384 37982 27396
rect 37976 27356 38021 27384
rect 37976 27344 37982 27356
rect 38286 27344 38292 27396
rect 38344 27384 38350 27396
rect 40221 27387 40279 27393
rect 38344 27356 39988 27384
rect 38344 27344 38350 27356
rect 28951 27288 29500 27316
rect 28951 27285 28963 27288
rect 28905 27279 28963 27285
rect 29546 27276 29552 27328
rect 29604 27316 29610 27328
rect 30101 27319 30159 27325
rect 30101 27316 30113 27319
rect 29604 27288 30113 27316
rect 29604 27276 29610 27288
rect 30101 27285 30113 27288
rect 30147 27285 30159 27319
rect 30101 27279 30159 27285
rect 30466 27276 30472 27328
rect 30524 27316 30530 27328
rect 30561 27319 30619 27325
rect 30561 27316 30573 27319
rect 30524 27288 30573 27316
rect 30524 27276 30530 27288
rect 30561 27285 30573 27288
rect 30607 27285 30619 27319
rect 31478 27316 31484 27328
rect 31439 27288 31484 27316
rect 30561 27279 30619 27285
rect 31478 27276 31484 27288
rect 31536 27276 31542 27328
rect 33962 27276 33968 27328
rect 34020 27316 34026 27328
rect 35802 27316 35808 27328
rect 34020 27288 35808 27316
rect 34020 27276 34026 27288
rect 35802 27276 35808 27288
rect 35860 27276 35866 27328
rect 38470 27316 38476 27328
rect 38431 27288 38476 27316
rect 38470 27276 38476 27288
rect 38528 27276 38534 27328
rect 38562 27276 38568 27328
rect 38620 27316 38626 27328
rect 39666 27316 39672 27328
rect 38620 27288 39672 27316
rect 38620 27276 38626 27288
rect 39666 27276 39672 27288
rect 39724 27276 39730 27328
rect 39850 27316 39856 27328
rect 39811 27288 39856 27316
rect 39850 27276 39856 27288
rect 39908 27276 39914 27328
rect 39960 27316 39988 27356
rect 40221 27353 40233 27387
rect 40267 27384 40279 27387
rect 40267 27356 40908 27384
rect 40267 27353 40279 27356
rect 40221 27347 40279 27353
rect 40880 27328 40908 27356
rect 41414 27344 41420 27396
rect 41472 27384 41478 27396
rect 46017 27387 46075 27393
rect 41472 27356 42748 27384
rect 41472 27344 41478 27356
rect 40313 27319 40371 27325
rect 40313 27316 40325 27319
rect 39960 27288 40325 27316
rect 40313 27285 40325 27288
rect 40359 27285 40371 27319
rect 40862 27316 40868 27328
rect 40823 27288 40868 27316
rect 40313 27279 40371 27285
rect 40862 27276 40868 27288
rect 40920 27276 40926 27328
rect 41141 27319 41199 27325
rect 41141 27285 41153 27319
rect 41187 27316 41199 27319
rect 41506 27316 41512 27328
rect 41187 27288 41512 27316
rect 41187 27285 41199 27288
rect 41141 27279 41199 27285
rect 41506 27276 41512 27288
rect 41564 27276 41570 27328
rect 41601 27319 41659 27325
rect 41601 27285 41613 27319
rect 41647 27316 41659 27319
rect 41966 27316 41972 27328
rect 41647 27288 41972 27316
rect 41647 27285 41659 27288
rect 41601 27279 41659 27285
rect 41966 27276 41972 27288
rect 42024 27276 42030 27328
rect 42610 27316 42616 27328
rect 42571 27288 42616 27316
rect 42610 27276 42616 27288
rect 42668 27276 42674 27328
rect 42720 27316 42748 27356
rect 46017 27353 46029 27387
rect 46063 27384 46075 27387
rect 46566 27384 46572 27396
rect 46063 27356 46572 27384
rect 46063 27353 46075 27356
rect 46017 27347 46075 27353
rect 46566 27344 46572 27356
rect 46624 27344 46630 27396
rect 46750 27344 46756 27396
rect 46808 27384 46814 27396
rect 49252 27384 49280 27424
rect 50154 27412 50160 27464
rect 50212 27452 50218 27464
rect 50525 27455 50583 27461
rect 50525 27452 50537 27455
rect 50212 27424 50537 27452
rect 50212 27412 50218 27424
rect 50525 27421 50537 27424
rect 50571 27421 50583 27455
rect 51169 27455 51227 27461
rect 51169 27452 51181 27455
rect 50525 27415 50583 27421
rect 50816 27424 51181 27452
rect 50614 27384 50620 27396
rect 46808 27356 49004 27384
rect 49252 27356 50620 27384
rect 46808 27344 46814 27356
rect 46109 27319 46167 27325
rect 46109 27316 46121 27319
rect 42720 27288 46121 27316
rect 46109 27285 46121 27288
rect 46155 27285 46167 27319
rect 46842 27316 46848 27328
rect 46803 27288 46848 27316
rect 46109 27279 46167 27285
rect 46842 27276 46848 27288
rect 46900 27276 46906 27328
rect 48222 27276 48228 27328
rect 48280 27316 48286 27328
rect 48774 27316 48780 27328
rect 48280 27288 48325 27316
rect 48735 27288 48780 27316
rect 48280 27276 48286 27288
rect 48774 27276 48780 27288
rect 48832 27276 48838 27328
rect 48976 27316 49004 27356
rect 50614 27344 50620 27356
rect 50672 27344 50678 27396
rect 50816 27384 50844 27424
rect 51169 27421 51181 27424
rect 51215 27421 51227 27455
rect 51169 27415 51227 27421
rect 52178 27412 52184 27464
rect 52236 27457 52242 27464
rect 52236 27412 52247 27457
rect 57149 27455 57207 27461
rect 57149 27421 57161 27455
rect 57195 27452 57207 27455
rect 57195 27424 57468 27452
rect 57195 27421 57207 27424
rect 57149 27415 57207 27421
rect 52189 27411 52247 27412
rect 50724 27356 50844 27384
rect 49145 27319 49203 27325
rect 49145 27316 49157 27319
rect 48976 27288 49157 27316
rect 49145 27285 49157 27288
rect 49191 27285 49203 27319
rect 49145 27279 49203 27285
rect 49237 27319 49295 27325
rect 49237 27285 49249 27319
rect 49283 27316 49295 27319
rect 50246 27316 50252 27328
rect 49283 27288 50252 27316
rect 49283 27285 49295 27288
rect 49237 27279 49295 27285
rect 50246 27276 50252 27288
rect 50304 27276 50310 27328
rect 50341 27319 50399 27325
rect 50341 27285 50353 27319
rect 50387 27316 50399 27319
rect 50724 27316 50752 27356
rect 54018 27344 54024 27396
rect 54076 27384 54082 27396
rect 54205 27387 54263 27393
rect 54205 27384 54217 27387
rect 54076 27356 54217 27384
rect 54076 27344 54082 27356
rect 54205 27353 54217 27356
rect 54251 27353 54263 27387
rect 54205 27347 54263 27353
rect 54941 27387 54999 27393
rect 54941 27353 54953 27387
rect 54987 27384 54999 27387
rect 54987 27356 55720 27384
rect 54987 27353 54999 27356
rect 54941 27347 54999 27353
rect 55692 27328 55720 27356
rect 57054 27344 57060 27396
rect 57112 27344 57118 27396
rect 57440 27384 57468 27424
rect 57698 27412 57704 27464
rect 57756 27452 57762 27464
rect 58158 27452 58164 27464
rect 57756 27424 58164 27452
rect 57756 27412 57762 27424
rect 58158 27412 58164 27424
rect 58216 27412 58222 27464
rect 58342 27452 58348 27464
rect 58303 27424 58348 27452
rect 58342 27412 58348 27424
rect 58400 27412 58406 27464
rect 58434 27412 58440 27464
rect 58492 27452 58498 27464
rect 58621 27455 58679 27461
rect 58621 27452 58633 27455
rect 58492 27424 58633 27452
rect 58492 27412 58498 27424
rect 58621 27421 58633 27424
rect 58667 27421 58679 27455
rect 58621 27415 58679 27421
rect 59354 27412 59360 27464
rect 59412 27452 59418 27464
rect 59817 27455 59875 27461
rect 59817 27452 59829 27455
rect 59412 27424 59829 27452
rect 59412 27412 59418 27424
rect 59817 27421 59829 27424
rect 59863 27421 59875 27455
rect 59817 27415 59875 27421
rect 60274 27412 60280 27464
rect 60332 27452 60338 27464
rect 60553 27455 60611 27461
rect 60553 27452 60565 27455
rect 60332 27424 60565 27452
rect 60332 27412 60338 27424
rect 60553 27421 60565 27424
rect 60599 27421 60611 27455
rect 60553 27415 60611 27421
rect 60829 27455 60887 27461
rect 60829 27421 60841 27455
rect 60875 27452 60887 27455
rect 61746 27452 61752 27464
rect 60875 27424 61752 27452
rect 60875 27421 60887 27424
rect 60829 27415 60887 27421
rect 61746 27412 61752 27424
rect 61804 27412 61810 27464
rect 62040 27461 62068 27492
rect 62114 27480 62120 27492
rect 62172 27480 62178 27532
rect 63218 27520 63224 27532
rect 63179 27492 63224 27520
rect 63218 27480 63224 27492
rect 63276 27480 63282 27532
rect 63310 27480 63316 27532
rect 63368 27520 63374 27532
rect 63368 27492 63632 27520
rect 63368 27480 63374 27492
rect 62025 27455 62083 27461
rect 62025 27421 62037 27455
rect 62071 27421 62083 27455
rect 63494 27452 63500 27464
rect 63455 27424 63500 27452
rect 62025 27415 62083 27421
rect 63494 27412 63500 27424
rect 63552 27412 63558 27464
rect 63604 27452 63632 27492
rect 64138 27480 64144 27532
rect 64196 27520 64202 27532
rect 64196 27492 65840 27520
rect 64196 27480 64202 27492
rect 64693 27455 64751 27461
rect 64693 27452 64705 27455
rect 63604 27424 64705 27452
rect 64693 27421 64705 27424
rect 64739 27421 64751 27455
rect 64693 27415 64751 27421
rect 64874 27412 64880 27464
rect 64932 27452 64938 27464
rect 65702 27452 65708 27464
rect 64932 27424 65708 27452
rect 64932 27412 64938 27424
rect 65702 27412 65708 27424
rect 65760 27412 65766 27464
rect 65812 27461 65840 27492
rect 68738 27480 68744 27532
rect 68796 27520 68802 27532
rect 68940 27520 68968 27560
rect 69014 27548 69020 27600
rect 69072 27588 69078 27600
rect 69385 27591 69443 27597
rect 69385 27588 69397 27591
rect 69072 27560 69397 27588
rect 69072 27548 69078 27560
rect 69385 27557 69397 27560
rect 69431 27557 69443 27591
rect 70486 27588 70492 27600
rect 69385 27551 69443 27557
rect 70136 27560 70492 27588
rect 70136 27520 70164 27560
rect 70486 27548 70492 27560
rect 70544 27548 70550 27600
rect 74626 27548 74632 27600
rect 74684 27588 74690 27600
rect 74684 27560 74729 27588
rect 74684 27548 74690 27560
rect 75270 27548 75276 27600
rect 75328 27588 75334 27600
rect 79778 27588 79784 27600
rect 75328 27560 79784 27588
rect 75328 27548 75334 27560
rect 79778 27548 79784 27560
rect 79836 27548 79842 27600
rect 81250 27548 81256 27600
rect 81308 27588 81314 27600
rect 81308 27560 81353 27588
rect 81308 27548 81314 27560
rect 81434 27548 81440 27600
rect 81492 27588 81498 27600
rect 81805 27591 81863 27597
rect 81805 27588 81817 27591
rect 81492 27560 81817 27588
rect 81492 27548 81498 27560
rect 81805 27557 81817 27560
rect 81851 27557 81863 27591
rect 82538 27588 82544 27600
rect 82499 27560 82544 27588
rect 81805 27551 81863 27557
rect 82538 27548 82544 27560
rect 82596 27548 82602 27600
rect 85574 27548 85580 27600
rect 85632 27588 85638 27600
rect 86221 27591 86279 27597
rect 86221 27588 86233 27591
rect 85632 27560 86233 27588
rect 85632 27548 85638 27560
rect 86221 27557 86233 27560
rect 86267 27557 86279 27591
rect 87046 27588 87052 27600
rect 87007 27560 87052 27588
rect 86221 27551 86279 27557
rect 87046 27548 87052 27560
rect 87104 27548 87110 27600
rect 87690 27588 87696 27600
rect 87651 27560 87696 27588
rect 87690 27548 87696 27560
rect 87748 27548 87754 27600
rect 95068 27588 95096 27628
rect 95896 27628 97304 27656
rect 101635 27628 101680 27656
rect 95786 27588 95792 27600
rect 89686 27560 95004 27588
rect 95068 27560 95792 27588
rect 68796 27492 68841 27520
rect 68940 27492 70164 27520
rect 68796 27480 68802 27492
rect 70394 27480 70400 27532
rect 70452 27520 70458 27532
rect 71317 27523 71375 27529
rect 71317 27520 71329 27523
rect 70452 27492 71329 27520
rect 70452 27480 70458 27492
rect 71317 27489 71329 27492
rect 71363 27489 71375 27523
rect 71317 27483 71375 27489
rect 71424 27492 72372 27520
rect 65797 27455 65855 27461
rect 65797 27421 65809 27455
rect 65843 27421 65855 27455
rect 65797 27415 65855 27421
rect 65886 27412 65892 27464
rect 65944 27452 65950 27464
rect 66441 27455 66499 27461
rect 66441 27452 66453 27455
rect 65944 27424 66453 27452
rect 65944 27412 65950 27424
rect 66441 27421 66453 27424
rect 66487 27421 66499 27455
rect 66441 27415 66499 27421
rect 66622 27412 66628 27464
rect 66680 27452 66686 27464
rect 67085 27455 67143 27461
rect 67085 27452 67097 27455
rect 66680 27424 67097 27452
rect 66680 27412 66686 27424
rect 67085 27421 67097 27424
rect 67131 27421 67143 27455
rect 67085 27415 67143 27421
rect 67821 27455 67879 27461
rect 67821 27421 67833 27455
rect 67867 27452 67879 27455
rect 68649 27455 68707 27461
rect 68649 27452 68661 27455
rect 67867 27424 68661 27452
rect 67867 27421 67879 27424
rect 67821 27415 67879 27421
rect 68649 27421 68661 27424
rect 68695 27452 68707 27455
rect 69290 27452 69296 27464
rect 68695 27424 69296 27452
rect 68695 27421 68707 27424
rect 68649 27415 68707 27421
rect 69290 27412 69296 27424
rect 69348 27412 69354 27464
rect 69474 27412 69480 27464
rect 69532 27452 69538 27464
rect 69569 27455 69627 27461
rect 69569 27452 69581 27455
rect 69532 27424 69581 27452
rect 69532 27412 69538 27424
rect 69569 27421 69581 27424
rect 69615 27421 69627 27455
rect 69569 27415 69627 27421
rect 70210 27412 70216 27464
rect 70268 27452 70274 27464
rect 71424 27452 71452 27492
rect 71958 27452 71964 27464
rect 70268 27424 70313 27452
rect 70504 27424 71452 27452
rect 71919 27424 71964 27452
rect 70268 27412 70274 27424
rect 58066 27384 58072 27396
rect 57440 27356 58072 27384
rect 58066 27344 58072 27356
rect 58124 27344 58130 27396
rect 59446 27384 59452 27396
rect 58360 27356 59452 27384
rect 50982 27316 50988 27328
rect 50387 27288 50752 27316
rect 50943 27288 50988 27316
rect 50387 27285 50399 27288
rect 50341 27279 50399 27285
rect 50982 27276 50988 27288
rect 51040 27276 51046 27328
rect 51902 27276 51908 27328
rect 51960 27316 51966 27328
rect 51997 27319 52055 27325
rect 51997 27316 52009 27319
rect 51960 27288 52009 27316
rect 51960 27276 51966 27288
rect 51997 27285 52009 27288
rect 52043 27285 52055 27319
rect 53190 27316 53196 27328
rect 53151 27288 53196 27316
rect 51997 27279 52055 27285
rect 53190 27276 53196 27288
rect 53248 27276 53254 27328
rect 53834 27316 53840 27328
rect 53795 27288 53840 27316
rect 53834 27276 53840 27288
rect 53892 27276 53898 27328
rect 55306 27276 55312 27328
rect 55364 27316 55370 27328
rect 55493 27319 55551 27325
rect 55493 27316 55505 27319
rect 55364 27288 55505 27316
rect 55364 27276 55370 27288
rect 55493 27285 55505 27288
rect 55539 27285 55551 27319
rect 55493 27279 55551 27285
rect 55674 27276 55680 27328
rect 55732 27316 55738 27328
rect 56410 27316 56416 27328
rect 55732 27288 56416 27316
rect 55732 27276 55738 27288
rect 56410 27276 56416 27288
rect 56468 27276 56474 27328
rect 57072 27316 57100 27344
rect 57241 27319 57299 27325
rect 57241 27316 57253 27319
rect 57072 27288 57253 27316
rect 57241 27285 57253 27288
rect 57287 27285 57299 27319
rect 57241 27279 57299 27285
rect 57606 27276 57612 27328
rect 57664 27316 57670 27328
rect 58360 27316 58388 27356
rect 59446 27344 59452 27356
rect 59504 27344 59510 27396
rect 59538 27344 59544 27396
rect 59596 27384 59602 27396
rect 59596 27356 59768 27384
rect 59596 27344 59602 27356
rect 57664 27288 58388 27316
rect 57664 27276 57670 27288
rect 59170 27276 59176 27328
rect 59228 27316 59234 27328
rect 59633 27319 59691 27325
rect 59633 27316 59645 27319
rect 59228 27288 59645 27316
rect 59228 27276 59234 27288
rect 59633 27285 59645 27288
rect 59679 27285 59691 27319
rect 59740 27316 59768 27356
rect 60642 27344 60648 27396
rect 60700 27384 60706 27396
rect 60700 27356 60964 27384
rect 60700 27344 60706 27356
rect 60826 27316 60832 27328
rect 59740 27288 60832 27316
rect 59633 27279 59691 27285
rect 60826 27276 60832 27288
rect 60884 27276 60890 27328
rect 60936 27316 60964 27356
rect 62040 27356 70256 27384
rect 62040 27316 62068 27356
rect 60936 27288 62068 27316
rect 62114 27276 62120 27328
rect 62172 27316 62178 27328
rect 64509 27319 64567 27325
rect 64509 27316 64521 27319
rect 62172 27288 64521 27316
rect 62172 27276 62178 27288
rect 64509 27285 64521 27288
rect 64555 27285 64567 27319
rect 64509 27279 64567 27285
rect 64598 27276 64604 27328
rect 64656 27316 64662 27328
rect 65613 27319 65671 27325
rect 65613 27316 65625 27319
rect 64656 27288 65625 27316
rect 64656 27276 64662 27288
rect 65613 27285 65625 27288
rect 65659 27285 65671 27319
rect 66254 27316 66260 27328
rect 66215 27288 66260 27316
rect 65613 27279 65671 27285
rect 66254 27276 66260 27288
rect 66312 27276 66318 27328
rect 66901 27319 66959 27325
rect 66901 27285 66913 27319
rect 66947 27316 66959 27319
rect 68002 27316 68008 27328
rect 66947 27288 68008 27316
rect 66947 27285 66959 27288
rect 66901 27279 66959 27285
rect 68002 27276 68008 27288
rect 68060 27276 68066 27328
rect 68186 27316 68192 27328
rect 68147 27288 68192 27316
rect 68186 27276 68192 27288
rect 68244 27276 68250 27328
rect 68462 27276 68468 27328
rect 68520 27316 68526 27328
rect 68557 27319 68615 27325
rect 68557 27316 68569 27319
rect 68520 27288 68569 27316
rect 68520 27276 68526 27288
rect 68557 27285 68569 27288
rect 68603 27285 68615 27319
rect 68557 27279 68615 27285
rect 69566 27276 69572 27328
rect 69624 27316 69630 27328
rect 70029 27319 70087 27325
rect 70029 27316 70041 27319
rect 69624 27288 70041 27316
rect 69624 27276 69630 27288
rect 70029 27285 70041 27288
rect 70075 27285 70087 27319
rect 70228 27316 70256 27356
rect 70504 27316 70532 27424
rect 71958 27412 71964 27424
rect 72016 27412 72022 27464
rect 72050 27412 72056 27464
rect 72108 27452 72114 27464
rect 72237 27455 72295 27461
rect 72237 27452 72249 27455
rect 72108 27424 72249 27452
rect 72108 27412 72114 27424
rect 72237 27421 72249 27424
rect 72283 27421 72295 27455
rect 72344 27452 72372 27492
rect 72418 27480 72424 27532
rect 72476 27520 72482 27532
rect 74902 27520 74908 27532
rect 72476 27492 74908 27520
rect 72476 27480 72482 27492
rect 74902 27480 74908 27492
rect 74960 27480 74966 27532
rect 75178 27520 75184 27532
rect 75139 27492 75184 27520
rect 75178 27480 75184 27492
rect 75236 27480 75242 27532
rect 75288 27492 77294 27520
rect 75288 27452 75316 27492
rect 72344 27424 75316 27452
rect 72237 27415 72295 27421
rect 75914 27412 75920 27464
rect 75972 27452 75978 27464
rect 76101 27455 76159 27461
rect 76101 27452 76113 27455
rect 75972 27424 76113 27452
rect 75972 27412 75978 27424
rect 76101 27421 76113 27424
rect 76147 27421 76159 27455
rect 76742 27452 76748 27464
rect 76703 27424 76748 27452
rect 76101 27415 76159 27421
rect 76742 27412 76748 27424
rect 76800 27412 76806 27464
rect 76834 27412 76840 27464
rect 76892 27452 76898 27464
rect 77021 27455 77079 27461
rect 77021 27452 77033 27455
rect 76892 27424 77033 27452
rect 76892 27412 76898 27424
rect 77021 27421 77033 27424
rect 77067 27421 77079 27455
rect 77266 27452 77294 27492
rect 78858 27480 78864 27532
rect 78916 27520 78922 27532
rect 79137 27523 79195 27529
rect 79137 27520 79149 27523
rect 78916 27492 79149 27520
rect 78916 27480 78922 27492
rect 79137 27489 79149 27492
rect 79183 27489 79195 27523
rect 79137 27483 79195 27489
rect 79321 27523 79379 27529
rect 79321 27489 79333 27523
rect 79367 27520 79379 27523
rect 79410 27520 79416 27532
rect 79367 27492 79416 27520
rect 79367 27489 79379 27492
rect 79321 27483 79379 27489
rect 79410 27480 79416 27492
rect 79468 27480 79474 27532
rect 84286 27480 84292 27532
rect 84344 27520 84350 27532
rect 85022 27520 85028 27532
rect 84344 27492 84884 27520
rect 84983 27492 85028 27520
rect 84344 27480 84350 27492
rect 77266 27424 79364 27452
rect 77021 27415 77079 27421
rect 70578 27344 70584 27396
rect 70636 27384 70642 27396
rect 78766 27384 78772 27396
rect 70636 27356 78772 27384
rect 70636 27344 70642 27356
rect 78766 27344 78772 27356
rect 78824 27344 78830 27396
rect 79336 27384 79364 27424
rect 79594 27412 79600 27464
rect 79652 27452 79658 27464
rect 80057 27455 80115 27461
rect 80057 27452 80069 27455
rect 79652 27424 80069 27452
rect 79652 27412 79658 27424
rect 80057 27421 80069 27424
rect 80103 27421 80115 27455
rect 80057 27415 80115 27421
rect 80514 27412 80520 27464
rect 80572 27452 80578 27464
rect 81069 27455 81127 27461
rect 81069 27452 81081 27455
rect 80572 27424 81081 27452
rect 80572 27412 80578 27424
rect 81069 27421 81081 27424
rect 81115 27421 81127 27455
rect 81986 27452 81992 27464
rect 81947 27424 81992 27452
rect 81069 27415 81127 27421
rect 81986 27412 81992 27424
rect 82044 27412 82050 27464
rect 82722 27452 82728 27464
rect 82683 27424 82728 27452
rect 82722 27412 82728 27424
rect 82780 27412 82786 27464
rect 83734 27412 83740 27464
rect 83792 27452 83798 27464
rect 83829 27455 83887 27461
rect 83829 27452 83841 27455
rect 83792 27424 83841 27452
rect 83792 27412 83798 27424
rect 83829 27421 83841 27424
rect 83875 27421 83887 27455
rect 83829 27415 83887 27421
rect 83918 27412 83924 27464
rect 83976 27452 83982 27464
rect 84856 27452 84884 27492
rect 85022 27480 85028 27492
rect 85080 27480 85086 27532
rect 85206 27480 85212 27532
rect 85264 27520 85270 27532
rect 89686 27520 89714 27560
rect 90634 27520 90640 27532
rect 85264 27492 89714 27520
rect 90595 27492 90640 27520
rect 85264 27480 85270 27492
rect 90634 27480 90640 27492
rect 90692 27480 90698 27532
rect 91370 27480 91376 27532
rect 91428 27520 91434 27532
rect 94866 27520 94872 27532
rect 91428 27492 94728 27520
rect 94827 27492 94872 27520
rect 91428 27480 91434 27492
rect 83976 27424 84792 27452
rect 84856 27424 86356 27452
rect 83976 27412 83982 27424
rect 84764 27384 84792 27424
rect 84841 27387 84899 27393
rect 84841 27384 84853 27387
rect 79336 27356 84608 27384
rect 84764 27356 84853 27384
rect 70228 27288 70532 27316
rect 70765 27319 70823 27325
rect 70029 27279 70087 27285
rect 70765 27285 70777 27319
rect 70811 27316 70823 27319
rect 70946 27316 70952 27328
rect 70811 27288 70952 27316
rect 70811 27285 70823 27288
rect 70765 27279 70823 27285
rect 70946 27276 70952 27288
rect 71004 27276 71010 27328
rect 71130 27316 71136 27328
rect 71091 27288 71136 27316
rect 71130 27276 71136 27288
rect 71188 27276 71194 27328
rect 71225 27319 71283 27325
rect 71225 27285 71237 27319
rect 71271 27316 71283 27319
rect 71314 27316 71320 27328
rect 71271 27288 71320 27316
rect 71271 27285 71283 27288
rect 71225 27279 71283 27285
rect 71314 27276 71320 27288
rect 71372 27276 71378 27328
rect 74258 27316 74264 27328
rect 74219 27288 74264 27316
rect 74258 27276 74264 27288
rect 74316 27316 74322 27328
rect 74534 27316 74540 27328
rect 74316 27288 74540 27316
rect 74316 27276 74322 27288
rect 74534 27276 74540 27288
rect 74592 27276 74598 27328
rect 74626 27276 74632 27328
rect 74684 27316 74690 27328
rect 74997 27319 75055 27325
rect 74997 27316 75009 27319
rect 74684 27288 75009 27316
rect 74684 27276 74690 27288
rect 74997 27285 75009 27288
rect 75043 27285 75055 27319
rect 74997 27279 75055 27285
rect 75089 27319 75147 27325
rect 75089 27285 75101 27319
rect 75135 27316 75147 27319
rect 75917 27319 75975 27325
rect 75917 27316 75929 27319
rect 75135 27288 75929 27316
rect 75135 27285 75147 27288
rect 75089 27279 75147 27285
rect 75917 27285 75929 27288
rect 75963 27285 75975 27319
rect 75917 27279 75975 27285
rect 76006 27276 76012 27328
rect 76064 27316 76070 27328
rect 78582 27316 78588 27328
rect 76064 27288 78588 27316
rect 76064 27276 76070 27288
rect 78582 27276 78588 27288
rect 78640 27276 78646 27328
rect 78677 27319 78735 27325
rect 78677 27285 78689 27319
rect 78723 27316 78735 27319
rect 78950 27316 78956 27328
rect 78723 27288 78956 27316
rect 78723 27285 78735 27288
rect 78677 27279 78735 27285
rect 78950 27276 78956 27288
rect 79008 27276 79014 27328
rect 79042 27276 79048 27328
rect 79100 27316 79106 27328
rect 79100 27288 79145 27316
rect 79100 27276 79106 27288
rect 79318 27276 79324 27328
rect 79376 27316 79382 27328
rect 79873 27319 79931 27325
rect 79873 27316 79885 27319
rect 79376 27288 79885 27316
rect 79376 27276 79382 27288
rect 79873 27285 79885 27288
rect 79919 27285 79931 27319
rect 79873 27279 79931 27285
rect 83645 27319 83703 27325
rect 83645 27285 83657 27319
rect 83691 27316 83703 27319
rect 84286 27316 84292 27328
rect 83691 27288 84292 27316
rect 83691 27285 83703 27288
rect 83645 27279 83703 27285
rect 84286 27276 84292 27288
rect 84344 27276 84350 27328
rect 84470 27316 84476 27328
rect 84431 27288 84476 27316
rect 84470 27276 84476 27288
rect 84528 27276 84534 27328
rect 84580 27316 84608 27356
rect 84841 27353 84853 27356
rect 84887 27353 84899 27387
rect 84841 27347 84899 27353
rect 84933 27387 84991 27393
rect 84933 27353 84945 27387
rect 84979 27384 84991 27387
rect 86126 27384 86132 27396
rect 84979 27356 86132 27384
rect 84979 27353 84991 27356
rect 84933 27347 84991 27353
rect 86126 27344 86132 27356
rect 86184 27344 86190 27396
rect 86328 27384 86356 27424
rect 86402 27412 86408 27464
rect 86460 27452 86466 27464
rect 87230 27452 87236 27464
rect 86460 27424 86505 27452
rect 87191 27424 87236 27452
rect 86460 27412 86466 27424
rect 87230 27412 87236 27424
rect 87288 27412 87294 27464
rect 87322 27412 87328 27464
rect 87380 27452 87386 27464
rect 87877 27455 87935 27461
rect 87877 27452 87889 27455
rect 87380 27424 87889 27452
rect 87380 27412 87386 27424
rect 87877 27421 87889 27424
rect 87923 27421 87935 27455
rect 87877 27415 87935 27421
rect 88334 27412 88340 27464
rect 88392 27452 88398 27464
rect 88981 27455 89039 27461
rect 88981 27452 88993 27455
rect 88392 27424 88993 27452
rect 88392 27412 88398 27424
rect 88981 27421 88993 27424
rect 89027 27421 89039 27455
rect 90545 27455 90603 27461
rect 90545 27452 90557 27455
rect 88981 27415 89039 27421
rect 90100 27424 90557 27452
rect 86954 27384 86960 27396
rect 86328 27356 86960 27384
rect 86954 27344 86960 27356
rect 87012 27344 87018 27396
rect 89349 27387 89407 27393
rect 89349 27384 89361 27387
rect 88628 27356 89361 27384
rect 88628 27316 88656 27356
rect 89349 27353 89361 27356
rect 89395 27353 89407 27387
rect 89349 27347 89407 27353
rect 88794 27316 88800 27328
rect 84580 27288 88656 27316
rect 88755 27288 88800 27316
rect 88794 27276 88800 27288
rect 88852 27276 88858 27328
rect 89364 27316 89392 27347
rect 89438 27344 89444 27396
rect 89496 27384 89502 27396
rect 89714 27384 89720 27396
rect 89496 27356 89720 27384
rect 89496 27344 89502 27356
rect 89714 27344 89720 27356
rect 89772 27344 89778 27396
rect 90100 27384 90128 27424
rect 90545 27421 90557 27424
rect 90591 27421 90603 27455
rect 90545 27415 90603 27421
rect 91462 27412 91468 27464
rect 91520 27452 91526 27464
rect 91833 27455 91891 27461
rect 91833 27452 91845 27455
rect 91520 27424 91845 27452
rect 91520 27412 91526 27424
rect 91833 27421 91845 27424
rect 91879 27421 91891 27455
rect 94590 27452 94596 27464
rect 91833 27415 91891 27421
rect 91940 27424 94596 27452
rect 91940 27384 91968 27424
rect 94590 27412 94596 27424
rect 94648 27412 94654 27464
rect 94700 27452 94728 27492
rect 94866 27480 94872 27492
rect 94924 27480 94930 27532
rect 94976 27520 95004 27560
rect 95786 27548 95792 27560
rect 95844 27548 95850 27600
rect 95896 27520 95924 27628
rect 95970 27548 95976 27600
rect 96028 27588 96034 27600
rect 96525 27591 96583 27597
rect 96525 27588 96537 27591
rect 96028 27560 96537 27588
rect 96028 27548 96034 27560
rect 96525 27557 96537 27560
rect 96571 27557 96583 27591
rect 96525 27551 96583 27557
rect 96890 27548 96896 27600
rect 96948 27588 96954 27600
rect 97169 27591 97227 27597
rect 97169 27588 97181 27591
rect 96948 27560 97181 27588
rect 96948 27548 96954 27560
rect 97169 27557 97181 27560
rect 97215 27557 97227 27591
rect 97169 27551 97227 27557
rect 94976 27492 95924 27520
rect 97276 27520 97304 27628
rect 101674 27616 101680 27628
rect 101732 27616 101738 27668
rect 97994 27588 98000 27600
rect 97955 27560 98000 27588
rect 97994 27548 98000 27560
rect 98052 27548 98058 27600
rect 98104 27560 99374 27588
rect 98104 27520 98132 27560
rect 97276 27492 98132 27520
rect 98546 27480 98552 27532
rect 98604 27520 98610 27532
rect 99101 27523 99159 27529
rect 99101 27520 99113 27523
rect 98604 27492 99113 27520
rect 98604 27480 98610 27492
rect 99101 27489 99113 27492
rect 99147 27489 99159 27523
rect 99346 27520 99374 27560
rect 99834 27548 99840 27600
rect 99892 27588 99898 27600
rect 100389 27591 100447 27597
rect 100389 27588 100401 27591
rect 99892 27560 100401 27588
rect 99892 27548 99898 27560
rect 100389 27557 100401 27560
rect 100435 27557 100447 27591
rect 100389 27551 100447 27557
rect 100938 27548 100944 27600
rect 100996 27588 101002 27600
rect 102505 27591 102563 27597
rect 102505 27588 102517 27591
rect 100996 27560 102517 27588
rect 100996 27548 101002 27560
rect 102505 27557 102517 27560
rect 102551 27557 102563 27591
rect 103146 27588 103152 27600
rect 103107 27560 103152 27588
rect 102505 27551 102563 27557
rect 103146 27548 103152 27560
rect 103204 27548 103210 27600
rect 105630 27548 105636 27600
rect 105688 27588 105694 27600
rect 106093 27591 106151 27597
rect 106093 27588 106105 27591
rect 105688 27560 106105 27588
rect 105688 27548 105694 27560
rect 106093 27557 106105 27560
rect 106139 27557 106151 27591
rect 106093 27551 106151 27557
rect 107654 27548 107660 27600
rect 107712 27588 107718 27600
rect 108301 27591 108359 27597
rect 108301 27588 108313 27591
rect 107712 27560 108313 27588
rect 107712 27548 107718 27560
rect 108301 27557 108313 27560
rect 108347 27557 108359 27591
rect 108301 27551 108359 27557
rect 109034 27548 109040 27600
rect 109092 27588 109098 27600
rect 109405 27591 109463 27597
rect 109405 27588 109417 27591
rect 109092 27560 109417 27588
rect 109092 27548 109098 27560
rect 109405 27557 109417 27560
rect 109451 27557 109463 27591
rect 109405 27551 109463 27557
rect 110877 27591 110935 27597
rect 110877 27557 110889 27591
rect 110923 27557 110935 27591
rect 113634 27588 113640 27600
rect 113595 27560 113640 27588
rect 110877 27551 110935 27557
rect 107473 27523 107531 27529
rect 107473 27520 107485 27523
rect 99346 27492 107485 27520
rect 99101 27483 99159 27489
rect 107473 27489 107485 27492
rect 107519 27520 107531 27523
rect 107749 27523 107807 27529
rect 107749 27520 107761 27523
rect 107519 27492 107761 27520
rect 107519 27489 107531 27492
rect 107473 27483 107531 27489
rect 107749 27489 107761 27492
rect 107795 27520 107807 27523
rect 108117 27523 108175 27529
rect 108117 27520 108129 27523
rect 107795 27492 108129 27520
rect 107795 27489 107807 27492
rect 107749 27483 107807 27489
rect 108117 27489 108129 27492
rect 108163 27489 108175 27523
rect 110892 27520 110920 27551
rect 113634 27548 113640 27560
rect 113692 27548 113698 27600
rect 115566 27588 115572 27600
rect 115527 27560 115572 27588
rect 115566 27548 115572 27560
rect 115624 27548 115630 27600
rect 108117 27483 108175 27489
rect 108224 27492 110920 27520
rect 95697 27455 95755 27461
rect 94700 27448 95648 27452
rect 95697 27448 95709 27455
rect 94700 27424 95709 27448
rect 95620 27421 95709 27424
rect 95743 27448 95755 27455
rect 95804 27448 96108 27452
rect 95743 27424 96108 27448
rect 95743 27421 95832 27424
rect 95620 27420 95832 27421
rect 95697 27415 95755 27420
rect 92750 27384 92756 27396
rect 89824 27356 90128 27384
rect 90376 27356 91968 27384
rect 92711 27356 92756 27384
rect 89824 27325 89852 27356
rect 89809 27319 89867 27325
rect 89809 27316 89821 27319
rect 89364 27288 89821 27316
rect 89809 27285 89821 27288
rect 89855 27285 89867 27319
rect 90082 27316 90088 27328
rect 90043 27288 90088 27316
rect 89809 27279 89867 27285
rect 90082 27276 90088 27288
rect 90140 27276 90146 27328
rect 90174 27276 90180 27328
rect 90232 27316 90238 27328
rect 90376 27316 90404 27356
rect 92750 27344 92756 27356
rect 92808 27344 92814 27396
rect 94777 27387 94835 27393
rect 94777 27353 94789 27387
rect 94823 27384 94835 27387
rect 96080 27384 96108 27424
rect 96706 27412 96712 27464
rect 96764 27452 96770 27464
rect 97353 27455 97411 27461
rect 97353 27452 97365 27455
rect 96764 27424 96809 27452
rect 96908 27424 97365 27452
rect 96764 27412 96770 27424
rect 94823 27356 96016 27384
rect 96080 27356 96384 27384
rect 94823 27353 94835 27356
rect 94777 27347 94835 27353
rect 90232 27288 90404 27316
rect 90453 27319 90511 27325
rect 90232 27276 90238 27288
rect 90453 27285 90465 27319
rect 90499 27316 90511 27319
rect 91002 27316 91008 27328
rect 90499 27288 91008 27316
rect 90499 27285 90511 27288
rect 90453 27279 90511 27285
rect 91002 27276 91008 27288
rect 91060 27276 91066 27328
rect 91922 27316 91928 27328
rect 91883 27288 91928 27316
rect 91922 27276 91928 27288
rect 91980 27276 91986 27328
rect 92842 27316 92848 27328
rect 92803 27288 92848 27316
rect 92842 27276 92848 27288
rect 92900 27276 92906 27328
rect 94317 27319 94375 27325
rect 94317 27285 94329 27319
rect 94363 27316 94375 27319
rect 94406 27316 94412 27328
rect 94363 27288 94412 27316
rect 94363 27285 94375 27288
rect 94317 27279 94375 27285
rect 94406 27276 94412 27288
rect 94464 27276 94470 27328
rect 94682 27316 94688 27328
rect 94643 27288 94688 27316
rect 94682 27276 94688 27288
rect 94740 27276 94746 27328
rect 94866 27276 94872 27328
rect 94924 27316 94930 27328
rect 95513 27319 95571 27325
rect 95513 27316 95525 27319
rect 94924 27288 95525 27316
rect 94924 27276 94930 27288
rect 95513 27285 95525 27288
rect 95559 27285 95571 27319
rect 95988 27316 96016 27356
rect 96246 27316 96252 27328
rect 95988 27288 96252 27316
rect 95513 27279 95571 27285
rect 96246 27276 96252 27288
rect 96304 27276 96310 27328
rect 96356 27316 96384 27356
rect 96430 27344 96436 27396
rect 96488 27384 96494 27396
rect 96908 27384 96936 27424
rect 97353 27421 97365 27424
rect 97399 27421 97411 27455
rect 98178 27452 98184 27464
rect 98139 27424 98184 27452
rect 97353 27415 97411 27421
rect 98178 27412 98184 27424
rect 98236 27412 98242 27464
rect 99374 27412 99380 27464
rect 99432 27452 99438 27464
rect 99432 27424 99477 27452
rect 99432 27412 99438 27424
rect 99558 27412 99564 27464
rect 99616 27452 99622 27464
rect 100573 27455 100631 27461
rect 100573 27452 100585 27455
rect 99616 27424 100585 27452
rect 99616 27412 99622 27424
rect 100573 27421 100585 27424
rect 100619 27421 100631 27455
rect 100573 27415 100631 27421
rect 101122 27412 101128 27464
rect 101180 27452 101186 27464
rect 101861 27455 101919 27461
rect 101861 27452 101873 27455
rect 101180 27424 101873 27452
rect 101180 27412 101186 27424
rect 101861 27421 101873 27424
rect 101907 27421 101919 27455
rect 102686 27452 102692 27464
rect 102647 27424 102692 27452
rect 101861 27415 101919 27421
rect 102686 27412 102692 27424
rect 102744 27412 102750 27464
rect 102778 27412 102784 27464
rect 102836 27452 102842 27464
rect 103333 27455 103391 27461
rect 103333 27452 103345 27455
rect 102836 27424 103345 27452
rect 102836 27412 102842 27424
rect 103333 27421 103345 27424
rect 103379 27421 103391 27455
rect 105354 27452 105360 27464
rect 105315 27424 105360 27452
rect 103333 27415 103391 27421
rect 105354 27412 105360 27424
rect 105412 27412 105418 27464
rect 106277 27455 106335 27461
rect 106277 27421 106289 27455
rect 106323 27452 106335 27455
rect 106366 27452 106372 27464
rect 106323 27424 106372 27452
rect 106323 27421 106335 27424
rect 106277 27415 106335 27421
rect 106366 27412 106372 27424
rect 106424 27412 106430 27464
rect 106918 27412 106924 27464
rect 106976 27452 106982 27464
rect 107289 27455 107347 27461
rect 107289 27452 107301 27455
rect 106976 27424 107301 27452
rect 106976 27412 106982 27424
rect 107289 27421 107301 27424
rect 107335 27421 107347 27455
rect 107289 27415 107347 27421
rect 96488 27356 96936 27384
rect 96488 27344 96494 27356
rect 97166 27344 97172 27396
rect 97224 27384 97230 27396
rect 100938 27384 100944 27396
rect 97224 27356 100944 27384
rect 97224 27344 97230 27356
rect 100938 27344 100944 27356
rect 100996 27344 101002 27396
rect 104710 27384 104716 27396
rect 104671 27356 104716 27384
rect 104710 27344 104716 27356
rect 104768 27344 104774 27396
rect 104986 27344 104992 27396
rect 105044 27384 105050 27396
rect 108224 27384 108252 27492
rect 110966 27480 110972 27532
rect 111024 27520 111030 27532
rect 116762 27520 116768 27532
rect 111024 27492 116768 27520
rect 111024 27480 111030 27492
rect 116762 27480 116768 27492
rect 116820 27480 116826 27532
rect 108482 27452 108488 27464
rect 108443 27424 108488 27452
rect 108482 27412 108488 27424
rect 108540 27412 108546 27464
rect 109586 27452 109592 27464
rect 109547 27424 109592 27452
rect 109586 27412 109592 27424
rect 109644 27412 109650 27464
rect 109770 27412 109776 27464
rect 109828 27452 109834 27464
rect 110233 27455 110291 27461
rect 110233 27452 110245 27455
rect 109828 27424 110245 27452
rect 109828 27412 109834 27424
rect 110233 27421 110245 27424
rect 110279 27421 110291 27455
rect 111058 27452 111064 27464
rect 111019 27424 111064 27452
rect 110233 27415 110291 27421
rect 111058 27412 111064 27424
rect 111116 27412 111122 27464
rect 112070 27412 112076 27464
rect 112128 27452 112134 27464
rect 112441 27455 112499 27461
rect 112441 27452 112453 27455
rect 112128 27424 112453 27452
rect 112128 27412 112134 27424
rect 112441 27421 112453 27424
rect 112487 27421 112499 27455
rect 112441 27415 112499 27421
rect 114554 27412 114560 27464
rect 114612 27452 114618 27464
rect 114741 27455 114799 27461
rect 114741 27452 114753 27455
rect 114612 27424 114753 27452
rect 114612 27412 114618 27424
rect 114741 27421 114753 27424
rect 114787 27421 114799 27455
rect 116026 27452 116032 27464
rect 115987 27424 116032 27452
rect 114741 27415 114799 27421
rect 116026 27412 116032 27424
rect 116084 27412 116090 27464
rect 117314 27452 117320 27464
rect 117275 27424 117320 27452
rect 117314 27412 117320 27424
rect 117372 27412 117378 27464
rect 117593 27455 117651 27461
rect 117593 27421 117605 27455
rect 117639 27421 117651 27455
rect 117593 27415 117651 27421
rect 117608 27384 117636 27415
rect 105044 27356 108252 27384
rect 109006 27356 117636 27384
rect 105044 27344 105050 27356
rect 96706 27316 96712 27328
rect 96356 27288 96712 27316
rect 96706 27276 96712 27288
rect 96764 27276 96770 27328
rect 104802 27316 104808 27328
rect 104763 27288 104808 27316
rect 104802 27276 104808 27288
rect 104860 27276 104866 27328
rect 104894 27276 104900 27328
rect 104952 27316 104958 27328
rect 105541 27319 105599 27325
rect 105541 27316 105553 27319
rect 104952 27288 105553 27316
rect 104952 27276 104958 27288
rect 105541 27285 105553 27288
rect 105587 27285 105599 27319
rect 105541 27279 105599 27285
rect 105630 27276 105636 27328
rect 105688 27316 105694 27328
rect 109006 27316 109034 27356
rect 110046 27316 110052 27328
rect 105688 27288 109034 27316
rect 110007 27288 110052 27316
rect 105688 27276 105694 27288
rect 110046 27276 110052 27288
rect 110104 27276 110110 27328
rect 112530 27316 112536 27328
rect 112491 27288 112536 27316
rect 112530 27276 112536 27288
rect 112588 27276 112594 27328
rect 114557 27319 114615 27325
rect 114557 27285 114569 27319
rect 114603 27316 114615 27319
rect 114738 27316 114744 27328
rect 114603 27288 114744 27316
rect 114603 27285 114615 27288
rect 114557 27279 114615 27285
rect 114738 27276 114744 27288
rect 114796 27276 114802 27328
rect 115198 27276 115204 27328
rect 115256 27316 115262 27328
rect 116213 27319 116271 27325
rect 116213 27316 116225 27319
rect 115256 27288 116225 27316
rect 115256 27276 115262 27288
rect 116213 27285 116225 27288
rect 116259 27285 116271 27319
rect 116213 27279 116271 27285
rect 1104 27226 118864 27248
rect 1104 27174 30398 27226
rect 30450 27174 30462 27226
rect 30514 27174 30526 27226
rect 30578 27174 30590 27226
rect 30642 27174 30654 27226
rect 30706 27174 59846 27226
rect 59898 27174 59910 27226
rect 59962 27174 59974 27226
rect 60026 27174 60038 27226
rect 60090 27174 60102 27226
rect 60154 27174 89294 27226
rect 89346 27174 89358 27226
rect 89410 27174 89422 27226
rect 89474 27174 89486 27226
rect 89538 27174 89550 27226
rect 89602 27174 118864 27226
rect 1104 27152 118864 27174
rect 1026 27072 1032 27124
rect 1084 27112 1090 27124
rect 3329 27115 3387 27121
rect 3329 27112 3341 27115
rect 1084 27084 3341 27112
rect 1084 27072 1090 27084
rect 3329 27081 3341 27084
rect 3375 27081 3387 27115
rect 4614 27112 4620 27124
rect 4575 27084 4620 27112
rect 3329 27075 3387 27081
rect 4614 27072 4620 27084
rect 4672 27072 4678 27124
rect 7834 27112 7840 27124
rect 7795 27084 7840 27112
rect 7834 27072 7840 27084
rect 7892 27072 7898 27124
rect 9674 27072 9680 27124
rect 9732 27112 9738 27124
rect 10597 27115 10655 27121
rect 10597 27112 10609 27115
rect 9732 27084 10609 27112
rect 9732 27072 9738 27084
rect 10597 27081 10609 27084
rect 10643 27081 10655 27115
rect 10597 27075 10655 27081
rect 11606 27072 11612 27124
rect 11664 27112 11670 27124
rect 11701 27115 11759 27121
rect 11701 27112 11713 27115
rect 11664 27084 11713 27112
rect 11664 27072 11670 27084
rect 11701 27081 11713 27084
rect 11747 27081 11759 27115
rect 26970 27112 26976 27124
rect 11701 27075 11759 27081
rect 11900 27084 26976 27112
rect 1302 26936 1308 26988
rect 1360 26976 1366 26988
rect 1397 26979 1455 26985
rect 1397 26976 1409 26979
rect 1360 26948 1409 26976
rect 1360 26936 1366 26948
rect 1397 26945 1409 26948
rect 1443 26945 1455 26979
rect 2866 26976 2872 26988
rect 2827 26948 2872 26976
rect 1397 26939 1455 26945
rect 2866 26936 2872 26948
rect 2924 26936 2930 26988
rect 3510 26976 3516 26988
rect 3471 26948 3516 26976
rect 3510 26936 3516 26948
rect 3568 26936 3574 26988
rect 4798 26976 4804 26988
rect 4759 26948 4804 26976
rect 4798 26936 4804 26948
rect 4856 26936 4862 26988
rect 8021 26979 8079 26985
rect 8021 26945 8033 26979
rect 8067 26945 8079 26979
rect 8021 26939 8079 26945
rect 1670 26908 1676 26920
rect 1631 26880 1676 26908
rect 1670 26868 1676 26880
rect 1728 26868 1734 26920
rect 8036 26908 8064 26939
rect 10226 26936 10232 26988
rect 10284 26976 10290 26988
rect 11900 26985 11928 27084
rect 26970 27072 26976 27084
rect 27028 27072 27034 27124
rect 27157 27115 27215 27121
rect 27157 27081 27169 27115
rect 27203 27112 27215 27115
rect 29178 27112 29184 27124
rect 27203 27084 29184 27112
rect 27203 27081 27215 27084
rect 27157 27075 27215 27081
rect 29178 27072 29184 27084
rect 29236 27072 29242 27124
rect 29365 27115 29423 27121
rect 29365 27081 29377 27115
rect 29411 27081 29423 27115
rect 29365 27075 29423 27081
rect 11974 27004 11980 27056
rect 12032 27044 12038 27056
rect 14458 27044 14464 27056
rect 12032 27016 14464 27044
rect 12032 27004 12038 27016
rect 14458 27004 14464 27016
rect 14516 27004 14522 27056
rect 15470 27004 15476 27056
rect 15528 27044 15534 27056
rect 15657 27047 15715 27053
rect 15657 27044 15669 27047
rect 15528 27016 15669 27044
rect 15528 27004 15534 27016
rect 15657 27013 15669 27016
rect 15703 27013 15715 27047
rect 15657 27007 15715 27013
rect 17126 27004 17132 27056
rect 17184 27044 17190 27056
rect 19702 27044 19708 27056
rect 17184 27016 19708 27044
rect 17184 27004 17190 27016
rect 19702 27004 19708 27016
rect 19760 27004 19766 27056
rect 22370 27004 22376 27056
rect 22428 27044 22434 27056
rect 26786 27044 26792 27056
rect 22428 27016 26792 27044
rect 22428 27004 22434 27016
rect 26786 27004 26792 27016
rect 26844 27004 26850 27056
rect 27062 27004 27068 27056
rect 27120 27044 27126 27056
rect 29270 27044 29276 27056
rect 27120 27016 29276 27044
rect 27120 27004 27126 27016
rect 29270 27004 29276 27016
rect 29328 27004 29334 27056
rect 10781 26979 10839 26985
rect 10781 26976 10793 26979
rect 10284 26948 10793 26976
rect 10284 26936 10290 26948
rect 10781 26945 10793 26948
rect 10827 26945 10839 26979
rect 10781 26939 10839 26945
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26945 11943 26979
rect 14274 26976 14280 26988
rect 14235 26948 14280 26976
rect 11885 26939 11943 26945
rect 14274 26936 14280 26948
rect 14332 26936 14338 26988
rect 14553 26979 14611 26985
rect 14553 26945 14565 26979
rect 14599 26976 14611 26979
rect 19794 26976 19800 26988
rect 14599 26948 19800 26976
rect 14599 26945 14611 26948
rect 14553 26939 14611 26945
rect 19794 26936 19800 26948
rect 19852 26936 19858 26988
rect 19889 26979 19947 26985
rect 19889 26945 19901 26979
rect 19935 26976 19947 26979
rect 20714 26976 20720 26988
rect 19935 26948 20720 26976
rect 19935 26945 19947 26948
rect 19889 26939 19947 26945
rect 20714 26936 20720 26948
rect 20772 26936 20778 26988
rect 27338 26976 27344 26988
rect 27299 26948 27344 26976
rect 27338 26936 27344 26948
rect 27396 26936 27402 26988
rect 29380 26976 29408 27075
rect 30466 27072 30472 27124
rect 30524 27112 30530 27124
rect 32674 27112 32680 27124
rect 30524 27084 32680 27112
rect 30524 27072 30530 27084
rect 32674 27072 32680 27084
rect 32732 27072 32738 27124
rect 32858 27072 32864 27124
rect 32916 27112 32922 27124
rect 32953 27115 33011 27121
rect 32953 27112 32965 27115
rect 32916 27084 32965 27112
rect 32916 27072 32922 27084
rect 32953 27081 32965 27084
rect 32999 27081 33011 27115
rect 33870 27112 33876 27124
rect 33831 27084 33876 27112
rect 32953 27075 33011 27081
rect 33870 27072 33876 27084
rect 33928 27072 33934 27124
rect 35253 27115 35311 27121
rect 35253 27112 35265 27115
rect 34072 27084 35265 27112
rect 31846 27004 31852 27056
rect 31904 27044 31910 27056
rect 33962 27044 33968 27056
rect 31904 27016 33968 27044
rect 31904 27004 31910 27016
rect 33962 27004 33968 27016
rect 34020 27004 34026 27056
rect 29546 26976 29552 26988
rect 27448 26948 29408 26976
rect 29507 26948 29552 26976
rect 24118 26908 24124 26920
rect 8036 26880 24124 26908
rect 24118 26868 24124 26880
rect 24176 26868 24182 26920
rect 27154 26868 27160 26920
rect 27212 26908 27218 26920
rect 27448 26908 27476 26948
rect 29546 26936 29552 26948
rect 29604 26936 29610 26988
rect 30377 26979 30435 26985
rect 30742 26980 30748 26988
rect 30377 26976 30389 26979
rect 29656 26948 30389 26976
rect 27212 26880 27476 26908
rect 27212 26868 27218 26880
rect 27522 26868 27528 26920
rect 27580 26908 27586 26920
rect 28994 26908 29000 26920
rect 27580 26880 29000 26908
rect 27580 26868 27586 26880
rect 28994 26868 29000 26880
rect 29052 26868 29058 26920
rect 29362 26868 29368 26920
rect 29420 26908 29426 26920
rect 29656 26908 29684 26948
rect 30377 26945 30389 26948
rect 30423 26945 30435 26979
rect 30668 26976 30748 26980
rect 30377 26939 30435 26945
rect 30576 26952 30748 26976
rect 30576 26948 30696 26952
rect 30576 26917 30604 26948
rect 30742 26936 30748 26952
rect 30800 26976 30806 26988
rect 32030 26976 32036 26988
rect 30800 26948 32036 26976
rect 30800 26936 30806 26948
rect 32030 26936 32036 26948
rect 32088 26936 32094 26988
rect 32122 26936 32128 26988
rect 32180 26976 32186 26988
rect 34072 26985 34100 27084
rect 35253 27081 35265 27084
rect 35299 27081 35311 27115
rect 35253 27075 35311 27081
rect 35434 27072 35440 27124
rect 35492 27112 35498 27124
rect 36449 27115 36507 27121
rect 36449 27112 36461 27115
rect 35492 27084 36461 27112
rect 35492 27072 35498 27084
rect 36449 27081 36461 27084
rect 36495 27081 36507 27115
rect 38102 27112 38108 27124
rect 38063 27084 38108 27112
rect 36449 27075 36507 27081
rect 38102 27072 38108 27084
rect 38160 27072 38166 27124
rect 38194 27072 38200 27124
rect 38252 27112 38258 27124
rect 40310 27112 40316 27124
rect 38252 27084 40316 27112
rect 38252 27072 38258 27084
rect 40310 27072 40316 27084
rect 40368 27072 40374 27124
rect 40494 27112 40500 27124
rect 40455 27084 40500 27112
rect 40494 27072 40500 27084
rect 40552 27072 40558 27124
rect 41322 27112 41328 27124
rect 41283 27084 41328 27112
rect 41322 27072 41328 27084
rect 41380 27072 41386 27124
rect 41598 27072 41604 27124
rect 41656 27112 41662 27124
rect 45646 27112 45652 27124
rect 41656 27084 45652 27112
rect 41656 27072 41662 27084
rect 45646 27072 45652 27084
rect 45704 27072 45710 27124
rect 45830 27112 45836 27124
rect 45791 27084 45836 27112
rect 45830 27072 45836 27084
rect 45888 27072 45894 27124
rect 52914 27112 52920 27124
rect 45940 27084 52776 27112
rect 52875 27084 52920 27112
rect 34882 27004 34888 27056
rect 34940 27044 34946 27056
rect 35621 27047 35679 27053
rect 35621 27044 35633 27047
rect 34940 27016 35633 27044
rect 34940 27004 34946 27016
rect 35621 27013 35633 27016
rect 35667 27013 35679 27047
rect 35621 27007 35679 27013
rect 38304 27016 41460 27044
rect 33137 26979 33195 26985
rect 33137 26976 33149 26979
rect 32180 26948 33149 26976
rect 32180 26936 32186 26948
rect 33137 26945 33149 26948
rect 33183 26945 33195 26979
rect 33137 26939 33195 26945
rect 34057 26979 34115 26985
rect 34057 26945 34069 26979
rect 34103 26945 34115 26979
rect 34606 26976 34612 26988
rect 34567 26948 34612 26976
rect 34057 26939 34115 26945
rect 34606 26936 34612 26948
rect 34664 26936 34670 26988
rect 35710 26976 35716 26988
rect 35671 26948 35716 26976
rect 35710 26936 35716 26948
rect 35768 26936 35774 26988
rect 35802 26936 35808 26988
rect 35860 26976 35866 26988
rect 36630 26976 36636 26988
rect 35860 26948 35940 26976
rect 36591 26948 36636 26976
rect 35860 26936 35866 26948
rect 35912 26917 35940 26948
rect 36630 26936 36636 26948
rect 36688 26936 36694 26988
rect 38304 26985 38332 27016
rect 41432 26988 41460 27016
rect 41874 27004 41880 27056
rect 41932 27044 41938 27056
rect 45940 27044 45968 27084
rect 46474 27044 46480 27056
rect 41932 27016 45968 27044
rect 46124 27016 46480 27044
rect 41932 27004 41938 27016
rect 38289 26979 38347 26985
rect 38289 26945 38301 26979
rect 38335 26945 38347 26979
rect 38289 26939 38347 26945
rect 38378 26936 38384 26988
rect 38436 26976 38442 26988
rect 38436 26948 39620 26976
rect 38436 26936 38442 26948
rect 30469 26911 30527 26917
rect 30469 26908 30481 26911
rect 29420 26880 29684 26908
rect 29748 26880 30481 26908
rect 29420 26868 29426 26880
rect 2685 26843 2743 26849
rect 2685 26809 2697 26843
rect 2731 26840 2743 26843
rect 2958 26840 2964 26852
rect 2731 26812 2964 26840
rect 2731 26809 2743 26812
rect 2685 26803 2743 26809
rect 2958 26800 2964 26812
rect 3016 26840 3022 26852
rect 9398 26840 9404 26852
rect 3016 26812 9404 26840
rect 3016 26800 3022 26812
rect 9398 26800 9404 26812
rect 9456 26800 9462 26852
rect 10502 26800 10508 26852
rect 10560 26840 10566 26852
rect 15841 26843 15899 26849
rect 10560 26812 15792 26840
rect 10560 26800 10566 26812
rect 9582 26732 9588 26784
rect 9640 26772 9646 26784
rect 15562 26772 15568 26784
rect 9640 26744 15568 26772
rect 9640 26732 9646 26744
rect 15562 26732 15568 26744
rect 15620 26732 15626 26784
rect 15764 26772 15792 26812
rect 15841 26809 15853 26843
rect 15887 26840 15899 26843
rect 16022 26840 16028 26852
rect 15887 26812 16028 26840
rect 15887 26809 15899 26812
rect 15841 26803 15899 26809
rect 16022 26800 16028 26812
rect 16080 26800 16086 26852
rect 17034 26800 17040 26852
rect 17092 26840 17098 26852
rect 20530 26840 20536 26852
rect 17092 26812 20116 26840
rect 20491 26812 20536 26840
rect 17092 26800 17098 26812
rect 19981 26775 20039 26781
rect 19981 26772 19993 26775
rect 15764 26744 19993 26772
rect 19981 26741 19993 26744
rect 20027 26741 20039 26775
rect 20088 26772 20116 26812
rect 20530 26800 20536 26812
rect 20588 26800 20594 26852
rect 22002 26800 22008 26852
rect 22060 26840 22066 26852
rect 22186 26840 22192 26852
rect 22060 26812 22192 26840
rect 22060 26800 22066 26812
rect 22186 26800 22192 26812
rect 22244 26800 22250 26852
rect 22278 26800 22284 26852
rect 22336 26840 22342 26852
rect 26786 26840 26792 26852
rect 22336 26812 26792 26840
rect 22336 26800 22342 26812
rect 26786 26800 26792 26812
rect 26844 26800 26850 26852
rect 27246 26800 27252 26852
rect 27304 26840 27310 26852
rect 29086 26840 29092 26852
rect 27304 26812 29092 26840
rect 27304 26800 27310 26812
rect 29086 26800 29092 26812
rect 29144 26800 29150 26852
rect 29546 26800 29552 26852
rect 29604 26840 29610 26852
rect 29748 26840 29776 26880
rect 30469 26877 30481 26880
rect 30515 26877 30527 26911
rect 30469 26871 30527 26877
rect 30561 26911 30619 26917
rect 30561 26877 30573 26911
rect 30607 26877 30619 26911
rect 35897 26911 35955 26917
rect 30561 26871 30619 26877
rect 33704 26880 34836 26908
rect 29604 26812 29776 26840
rect 30009 26843 30067 26849
rect 29604 26800 29610 26812
rect 30009 26809 30021 26843
rect 30055 26840 30067 26843
rect 33594 26840 33600 26852
rect 30055 26812 33600 26840
rect 30055 26809 30067 26812
rect 30009 26803 30067 26809
rect 33594 26800 33600 26812
rect 33652 26800 33658 26852
rect 21082 26772 21088 26784
rect 20088 26744 21088 26772
rect 19981 26735 20039 26741
rect 21082 26732 21088 26744
rect 21140 26732 21146 26784
rect 21910 26732 21916 26784
rect 21968 26772 21974 26784
rect 27062 26772 27068 26784
rect 21968 26744 27068 26772
rect 21968 26732 21974 26744
rect 27062 26732 27068 26744
rect 27120 26732 27126 26784
rect 27154 26732 27160 26784
rect 27212 26772 27218 26784
rect 29270 26772 29276 26784
rect 27212 26744 29276 26772
rect 27212 26732 27218 26744
rect 29270 26732 29276 26744
rect 29328 26732 29334 26784
rect 30098 26732 30104 26784
rect 30156 26772 30162 26784
rect 33704 26772 33732 26880
rect 30156 26744 33732 26772
rect 30156 26732 30162 26744
rect 34054 26732 34060 26784
rect 34112 26772 34118 26784
rect 34701 26775 34759 26781
rect 34701 26772 34713 26775
rect 34112 26744 34713 26772
rect 34112 26732 34118 26744
rect 34701 26741 34713 26744
rect 34747 26741 34759 26775
rect 34808 26772 34836 26880
rect 35897 26877 35909 26911
rect 35943 26877 35955 26911
rect 35897 26871 35955 26877
rect 39209 26911 39267 26917
rect 39209 26877 39221 26911
rect 39255 26877 39267 26911
rect 39209 26871 39267 26877
rect 34974 26800 34980 26852
rect 35032 26840 35038 26852
rect 39224 26840 39252 26871
rect 39298 26868 39304 26920
rect 39356 26908 39362 26920
rect 39485 26911 39543 26917
rect 39485 26908 39497 26911
rect 39356 26880 39497 26908
rect 39356 26868 39362 26880
rect 39485 26877 39497 26880
rect 39531 26877 39543 26911
rect 39485 26871 39543 26877
rect 35032 26812 39252 26840
rect 39592 26840 39620 26948
rect 39850 26936 39856 26988
rect 39908 26976 39914 26988
rect 40681 26979 40739 26985
rect 40681 26976 40693 26979
rect 39908 26948 40693 26976
rect 39908 26936 39914 26948
rect 40681 26945 40693 26948
rect 40727 26945 40739 26979
rect 40681 26939 40739 26945
rect 41414 26936 41420 26988
rect 41472 26936 41478 26988
rect 41509 26983 41567 26989
rect 41509 26949 41521 26983
rect 41555 26949 41567 26983
rect 41509 26943 41567 26949
rect 46017 26979 46075 26985
rect 46017 26945 46029 26979
rect 46063 26976 46075 26979
rect 46124 26976 46152 27016
rect 46474 27004 46480 27016
rect 46532 27004 46538 27056
rect 46566 27004 46572 27056
rect 46624 27044 46630 27056
rect 46661 27047 46719 27053
rect 46661 27044 46673 27047
rect 46624 27016 46673 27044
rect 46624 27004 46630 27016
rect 46661 27013 46673 27016
rect 46707 27013 46719 27047
rect 46661 27007 46719 27013
rect 46842 27004 46848 27056
rect 46900 27044 46906 27056
rect 50614 27044 50620 27056
rect 46900 27016 50620 27044
rect 46900 27004 46906 27016
rect 50614 27004 50620 27016
rect 50672 27004 50678 27056
rect 50706 27004 50712 27056
rect 50764 27044 50770 27056
rect 50764 27016 50809 27044
rect 50764 27004 50770 27016
rect 51166 27004 51172 27056
rect 51224 27004 51230 27056
rect 46063 26948 46152 26976
rect 46063 26945 46075 26948
rect 39666 26868 39672 26920
rect 39724 26908 39730 26920
rect 41230 26908 41236 26920
rect 39724 26880 41236 26908
rect 39724 26868 39730 26880
rect 41230 26868 41236 26880
rect 41288 26868 41294 26920
rect 41524 26908 41552 26943
rect 46017 26939 46075 26945
rect 46198 26936 46204 26988
rect 46256 26976 46262 26988
rect 46256 26948 48912 26976
rect 46256 26936 46262 26948
rect 41690 26908 41696 26920
rect 41524 26880 41696 26908
rect 41690 26868 41696 26880
rect 41748 26868 41754 26920
rect 48041 26911 48099 26917
rect 48041 26908 48053 26911
rect 41800 26880 48053 26908
rect 41800 26840 41828 26880
rect 48041 26877 48053 26880
rect 48087 26877 48099 26911
rect 48041 26871 48099 26877
rect 48317 26911 48375 26917
rect 48317 26877 48329 26911
rect 48363 26908 48375 26911
rect 48498 26908 48504 26920
rect 48363 26880 48504 26908
rect 48363 26877 48375 26880
rect 48317 26871 48375 26877
rect 48498 26868 48504 26880
rect 48556 26868 48562 26920
rect 48884 26908 48912 26948
rect 48958 26936 48964 26988
rect 49016 26976 49022 26988
rect 49513 26979 49571 26985
rect 49513 26976 49525 26979
rect 49016 26948 49525 26976
rect 49016 26936 49022 26948
rect 49513 26945 49525 26948
rect 49559 26945 49571 26979
rect 49513 26939 49571 26945
rect 50062 26936 50068 26988
rect 50120 26976 50126 26988
rect 50157 26979 50215 26985
rect 50157 26976 50169 26979
rect 50120 26948 50169 26976
rect 50120 26936 50126 26948
rect 50157 26945 50169 26948
rect 50203 26945 50215 26979
rect 50157 26939 50215 26945
rect 50338 26936 50344 26988
rect 50396 26976 50402 26988
rect 50724 26976 50752 27004
rect 50396 26948 50752 26976
rect 50893 26979 50951 26985
rect 50396 26936 50402 26948
rect 50893 26945 50905 26979
rect 50939 26976 50951 26979
rect 51184 26976 51212 27004
rect 50939 26948 51212 26976
rect 51445 26979 51503 26985
rect 50939 26945 50951 26948
rect 50893 26939 50951 26945
rect 51445 26945 51457 26979
rect 51491 26945 51503 26979
rect 51445 26939 51503 26945
rect 50706 26908 50712 26920
rect 48884 26880 50712 26908
rect 50706 26868 50712 26880
rect 50764 26868 50770 26920
rect 51460 26908 51488 26939
rect 50816 26880 51488 26908
rect 51629 26911 51687 26917
rect 39592 26812 41828 26840
rect 35032 26800 35038 26812
rect 44082 26800 44088 26852
rect 44140 26840 44146 26852
rect 45922 26840 45928 26852
rect 44140 26812 45928 26840
rect 44140 26800 44146 26812
rect 45922 26800 45928 26812
rect 45980 26800 45986 26852
rect 49970 26840 49976 26852
rect 46032 26812 49832 26840
rect 49931 26812 49976 26840
rect 46032 26772 46060 26812
rect 46934 26772 46940 26784
rect 34808 26744 46060 26772
rect 46895 26744 46940 26772
rect 34701 26735 34759 26741
rect 46934 26732 46940 26744
rect 46992 26732 46998 26784
rect 47118 26732 47124 26784
rect 47176 26772 47182 26784
rect 49050 26772 49056 26784
rect 47176 26744 49056 26772
rect 47176 26732 47182 26744
rect 49050 26732 49056 26744
rect 49108 26732 49114 26784
rect 49142 26732 49148 26784
rect 49200 26772 49206 26784
rect 49329 26775 49387 26781
rect 49329 26772 49341 26775
rect 49200 26744 49341 26772
rect 49200 26732 49206 26744
rect 49329 26741 49341 26744
rect 49375 26741 49387 26775
rect 49804 26772 49832 26812
rect 49970 26800 49976 26812
rect 50028 26800 50034 26852
rect 50154 26800 50160 26852
rect 50212 26840 50218 26852
rect 50816 26840 50844 26880
rect 51629 26877 51641 26911
rect 51675 26908 51687 26911
rect 51718 26908 51724 26920
rect 51675 26880 51724 26908
rect 51675 26877 51687 26880
rect 51629 26871 51687 26877
rect 51718 26868 51724 26880
rect 51776 26868 51782 26920
rect 52748 26908 52776 27084
rect 52914 27072 52920 27084
rect 52972 27072 52978 27124
rect 53006 27072 53012 27124
rect 53064 27112 53070 27124
rect 53064 27084 53972 27112
rect 53064 27072 53070 27084
rect 53282 27044 53288 27056
rect 53116 27016 53288 27044
rect 53116 26985 53144 27016
rect 53282 27004 53288 27016
rect 53340 27004 53346 27056
rect 53377 27047 53435 27053
rect 53377 27013 53389 27047
rect 53423 27044 53435 27047
rect 53834 27044 53840 27056
rect 53423 27016 53840 27044
rect 53423 27013 53435 27016
rect 53377 27007 53435 27013
rect 53834 27004 53840 27016
rect 53892 27004 53898 27056
rect 53944 27044 53972 27084
rect 54018 27072 54024 27124
rect 54076 27112 54082 27124
rect 55309 27115 55367 27121
rect 55309 27112 55321 27115
rect 54076 27084 55321 27112
rect 54076 27072 54082 27084
rect 55309 27081 55321 27084
rect 55355 27081 55367 27115
rect 55309 27075 55367 27081
rect 55398 27072 55404 27124
rect 55456 27112 55462 27124
rect 56137 27115 56195 27121
rect 56137 27112 56149 27115
rect 55456 27084 56149 27112
rect 55456 27072 55462 27084
rect 56137 27081 56149 27084
rect 56183 27081 56195 27115
rect 56502 27112 56508 27124
rect 56463 27084 56508 27112
rect 56137 27075 56195 27081
rect 56502 27072 56508 27084
rect 56560 27072 56566 27124
rect 57149 27115 57207 27121
rect 57149 27081 57161 27115
rect 57195 27112 57207 27115
rect 57514 27112 57520 27124
rect 57195 27084 57520 27112
rect 57195 27081 57207 27084
rect 57149 27075 57207 27081
rect 57514 27072 57520 27084
rect 57572 27072 57578 27124
rect 58066 27072 58072 27124
rect 58124 27112 58130 27124
rect 58345 27115 58403 27121
rect 58345 27112 58357 27115
rect 58124 27084 58357 27112
rect 58124 27072 58130 27084
rect 58345 27081 58357 27084
rect 58391 27081 58403 27115
rect 58345 27075 58403 27081
rect 58526 27072 58532 27124
rect 58584 27112 58590 27124
rect 58805 27115 58863 27121
rect 58805 27112 58817 27115
rect 58584 27084 58817 27112
rect 58584 27072 58590 27084
rect 58805 27081 58817 27084
rect 58851 27081 58863 27115
rect 59170 27112 59176 27124
rect 59131 27084 59176 27112
rect 58805 27075 58863 27081
rect 59170 27072 59176 27084
rect 59228 27072 59234 27124
rect 70486 27112 70492 27124
rect 62592 27084 70492 27112
rect 59078 27044 59084 27056
rect 53944 27016 59084 27044
rect 59078 27004 59084 27016
rect 59136 27004 59142 27056
rect 59446 27004 59452 27056
rect 59504 27044 59510 27056
rect 62592 27044 62620 27084
rect 70486 27072 70492 27084
rect 70544 27072 70550 27124
rect 71130 27072 71136 27124
rect 71188 27112 71194 27124
rect 74534 27112 74540 27124
rect 71188 27084 74540 27112
rect 71188 27072 71194 27084
rect 74534 27072 74540 27084
rect 74592 27072 74598 27124
rect 74718 27072 74724 27124
rect 74776 27112 74782 27124
rect 77021 27115 77079 27121
rect 74776 27084 76144 27112
rect 74776 27072 74782 27084
rect 59504 27016 62620 27044
rect 59504 27004 59510 27016
rect 62942 27004 62948 27056
rect 63000 27044 63006 27056
rect 64877 27047 64935 27053
rect 64877 27044 64889 27047
rect 63000 27016 64889 27044
rect 63000 27004 63006 27016
rect 64877 27013 64889 27016
rect 64923 27013 64935 27047
rect 64877 27007 64935 27013
rect 64984 27016 66668 27044
rect 53101 26979 53159 26985
rect 53101 26945 53113 26979
rect 53147 26945 53159 26979
rect 53101 26939 53159 26945
rect 53208 26948 54156 26976
rect 53208 26908 53236 26948
rect 52748 26880 53236 26908
rect 53653 26911 53711 26917
rect 53653 26877 53665 26911
rect 53699 26877 53711 26911
rect 53926 26908 53932 26920
rect 53887 26880 53932 26908
rect 53653 26871 53711 26877
rect 53668 26840 53696 26871
rect 53926 26868 53932 26880
rect 53984 26868 53990 26920
rect 54018 26840 54024 26852
rect 50212 26812 50844 26840
rect 51046 26812 53604 26840
rect 53668 26812 54024 26840
rect 50212 26800 50218 26812
rect 51046 26772 51074 26812
rect 49804 26744 51074 26772
rect 49329 26735 49387 26741
rect 51626 26732 51632 26784
rect 51684 26772 51690 26784
rect 53469 26775 53527 26781
rect 53469 26772 53481 26775
rect 51684 26744 53481 26772
rect 51684 26732 51690 26744
rect 53469 26741 53481 26744
rect 53515 26741 53527 26775
rect 53576 26772 53604 26812
rect 54018 26800 54024 26812
rect 54076 26800 54082 26852
rect 54128 26840 54156 26948
rect 55122 26936 55128 26988
rect 55180 26976 55186 26988
rect 55490 26976 55496 26988
rect 55180 26948 55496 26976
rect 55180 26936 55186 26948
rect 55490 26936 55496 26948
rect 55548 26936 55554 26988
rect 55674 26976 55680 26988
rect 55635 26948 55680 26976
rect 55674 26936 55680 26948
rect 55732 26936 55738 26988
rect 56318 26976 56324 26988
rect 56279 26948 56324 26976
rect 56318 26936 56324 26948
rect 56376 26936 56382 26988
rect 56686 26976 56692 26988
rect 56647 26948 56692 26976
rect 56686 26936 56692 26948
rect 56744 26936 56750 26988
rect 57330 26976 57336 26988
rect 57291 26948 57336 26976
rect 57330 26936 57336 26948
rect 57388 26936 57394 26988
rect 59170 26976 59176 26988
rect 57440 26948 59176 26976
rect 54294 26868 54300 26920
rect 54352 26908 54358 26920
rect 55769 26911 55827 26917
rect 55769 26908 55781 26911
rect 54352 26880 55781 26908
rect 54352 26868 54358 26880
rect 55769 26877 55781 26880
rect 55815 26877 55827 26911
rect 55769 26871 55827 26877
rect 55858 26868 55864 26920
rect 55916 26908 55922 26920
rect 57238 26908 57244 26920
rect 55916 26880 57244 26908
rect 55916 26868 55922 26880
rect 57238 26868 57244 26880
rect 57296 26868 57302 26920
rect 57440 26840 57468 26948
rect 59170 26936 59176 26948
rect 59228 26936 59234 26988
rect 59265 26979 59323 26985
rect 59265 26945 59277 26979
rect 59311 26976 59323 26979
rect 59354 26976 59360 26988
rect 59311 26948 59360 26976
rect 59311 26945 59323 26948
rect 59265 26939 59323 26945
rect 59354 26936 59360 26948
rect 59412 26936 59418 26988
rect 59630 26976 59636 26988
rect 59464 26948 59636 26976
rect 57885 26911 57943 26917
rect 57885 26877 57897 26911
rect 57931 26908 57943 26911
rect 58066 26908 58072 26920
rect 57931 26880 58072 26908
rect 57931 26877 57943 26880
rect 57885 26871 57943 26877
rect 58066 26868 58072 26880
rect 58124 26868 58130 26920
rect 58250 26868 58256 26920
rect 58308 26908 58314 26920
rect 59464 26917 59492 26948
rect 59630 26936 59636 26948
rect 59688 26936 59694 26988
rect 60001 26979 60059 26985
rect 60001 26945 60013 26979
rect 60047 26976 60059 26979
rect 60182 26976 60188 26988
rect 60047 26948 60188 26976
rect 60047 26945 60059 26948
rect 60001 26939 60059 26945
rect 60182 26936 60188 26948
rect 60240 26936 60246 26988
rect 61746 26976 61752 26988
rect 60384 26948 61752 26976
rect 59449 26911 59507 26917
rect 58308 26880 58388 26908
rect 58308 26868 58314 26880
rect 58158 26840 58164 26852
rect 54128 26812 57468 26840
rect 58119 26812 58164 26840
rect 58158 26800 58164 26812
rect 58216 26800 58222 26852
rect 58360 26840 58388 26880
rect 59449 26877 59461 26911
rect 59495 26877 59507 26911
rect 59449 26871 59507 26877
rect 59538 26868 59544 26920
rect 59596 26908 59602 26920
rect 60277 26911 60335 26917
rect 60277 26908 60289 26911
rect 59596 26880 60289 26908
rect 59596 26868 59602 26880
rect 60277 26877 60289 26880
rect 60323 26877 60335 26911
rect 60277 26871 60335 26877
rect 60384 26840 60412 26948
rect 61746 26936 61752 26948
rect 61804 26936 61810 26988
rect 61930 26976 61936 26988
rect 61891 26948 61936 26976
rect 61930 26936 61936 26948
rect 61988 26936 61994 26988
rect 62574 26976 62580 26988
rect 62535 26948 62580 26976
rect 62574 26936 62580 26948
rect 62632 26976 62638 26988
rect 62776 26976 62896 26980
rect 63678 26976 63684 26988
rect 62632 26952 63684 26976
rect 62632 26948 62804 26952
rect 62868 26948 63684 26952
rect 62632 26936 62638 26948
rect 63678 26936 63684 26948
rect 63736 26936 63742 26988
rect 63773 26979 63831 26985
rect 63773 26945 63785 26979
rect 63819 26976 63831 26979
rect 64598 26976 64604 26988
rect 63819 26948 64604 26976
rect 63819 26945 63831 26948
rect 63773 26939 63831 26945
rect 64598 26936 64604 26948
rect 64656 26936 64662 26988
rect 64690 26936 64696 26988
rect 64748 26976 64754 26988
rect 64984 26976 65012 27016
rect 65889 26979 65947 26985
rect 65889 26976 65901 26979
rect 64748 26948 65012 26976
rect 65260 26948 65901 26976
rect 64748 26936 64754 26948
rect 60458 26868 60464 26920
rect 60516 26908 60522 26920
rect 62025 26911 62083 26917
rect 62025 26908 62037 26911
rect 60516 26880 62037 26908
rect 60516 26868 60522 26880
rect 62025 26877 62037 26880
rect 62071 26877 62083 26911
rect 62206 26908 62212 26920
rect 62167 26880 62212 26908
rect 62025 26871 62083 26877
rect 62206 26868 62212 26880
rect 62264 26868 62270 26920
rect 62390 26868 62396 26920
rect 62448 26908 62454 26920
rect 63865 26911 63923 26917
rect 63865 26908 63877 26911
rect 62448 26880 63877 26908
rect 62448 26868 62454 26880
rect 63865 26877 63877 26880
rect 63911 26908 63923 26911
rect 63911 26880 64828 26908
rect 63911 26877 63923 26880
rect 63865 26871 63923 26877
rect 58360 26812 60412 26840
rect 60550 26800 60556 26852
rect 60608 26840 60614 26852
rect 60608 26812 60964 26840
rect 60608 26800 60614 26812
rect 54294 26772 54300 26784
rect 53576 26744 54300 26772
rect 53469 26735 53527 26741
rect 54294 26732 54300 26744
rect 54352 26732 54358 26784
rect 54386 26732 54392 26784
rect 54444 26772 54450 26784
rect 60642 26772 60648 26784
rect 54444 26744 60648 26772
rect 54444 26732 54450 26744
rect 60642 26732 60648 26744
rect 60700 26732 60706 26784
rect 60936 26772 60964 26812
rect 61194 26800 61200 26852
rect 61252 26840 61258 26852
rect 64690 26840 64696 26852
rect 61252 26812 64696 26840
rect 61252 26800 61258 26812
rect 64690 26800 64696 26812
rect 64748 26800 64754 26852
rect 64800 26840 64828 26880
rect 64874 26868 64880 26920
rect 64932 26908 64938 26920
rect 64969 26911 65027 26917
rect 64969 26908 64981 26911
rect 64932 26880 64981 26908
rect 64932 26868 64938 26880
rect 64969 26877 64981 26880
rect 65015 26877 65027 26911
rect 64969 26871 65027 26877
rect 65061 26911 65119 26917
rect 65061 26877 65073 26911
rect 65107 26877 65119 26911
rect 65061 26871 65119 26877
rect 65076 26840 65104 26871
rect 64800 26812 65104 26840
rect 61470 26772 61476 26784
rect 60936 26744 61476 26772
rect 61470 26732 61476 26744
rect 61528 26732 61534 26784
rect 61565 26775 61623 26781
rect 61565 26741 61577 26775
rect 61611 26772 61623 26775
rect 61838 26772 61844 26784
rect 61611 26744 61844 26772
rect 61611 26741 61623 26744
rect 61565 26735 61623 26741
rect 61838 26732 61844 26744
rect 61896 26732 61902 26784
rect 61930 26732 61936 26784
rect 61988 26772 61994 26784
rect 63218 26772 63224 26784
rect 61988 26744 63224 26772
rect 61988 26732 61994 26744
rect 63218 26732 63224 26744
rect 63276 26732 63282 26784
rect 63313 26775 63371 26781
rect 63313 26741 63325 26775
rect 63359 26772 63371 26775
rect 64046 26772 64052 26784
rect 63359 26744 64052 26772
rect 63359 26741 63371 26744
rect 63313 26735 63371 26741
rect 64046 26732 64052 26744
rect 64104 26732 64110 26784
rect 64138 26732 64144 26784
rect 64196 26772 64202 26784
rect 64325 26775 64383 26781
rect 64325 26772 64337 26775
rect 64196 26744 64337 26772
rect 64196 26732 64202 26744
rect 64325 26741 64337 26744
rect 64371 26741 64383 26775
rect 64325 26735 64383 26741
rect 64509 26775 64567 26781
rect 64509 26741 64521 26775
rect 64555 26772 64567 26775
rect 65260 26772 65288 26948
rect 65889 26945 65901 26948
rect 65935 26945 65947 26979
rect 65889 26939 65947 26945
rect 65978 26936 65984 26988
rect 66036 26976 66042 26988
rect 66533 26979 66591 26985
rect 66533 26976 66545 26979
rect 66036 26948 66545 26976
rect 66036 26936 66042 26948
rect 66533 26945 66545 26948
rect 66579 26945 66591 26979
rect 66640 26976 66668 27016
rect 68186 27004 68192 27056
rect 68244 27044 68250 27056
rect 68649 27047 68707 27053
rect 68649 27044 68661 27047
rect 68244 27016 68661 27044
rect 68244 27004 68250 27016
rect 68649 27013 68661 27016
rect 68695 27013 68707 27047
rect 70305 27047 70363 27053
rect 70305 27044 70317 27047
rect 68649 27007 68707 27013
rect 68756 27016 70317 27044
rect 68756 26976 68784 27016
rect 70305 27013 70317 27016
rect 70351 27013 70363 27047
rect 70305 27007 70363 27013
rect 71866 27004 71872 27056
rect 71924 27044 71930 27056
rect 71924 27016 72740 27044
rect 71924 27004 71930 27016
rect 66640 26948 68784 26976
rect 66533 26939 66591 26945
rect 68830 26936 68836 26988
rect 68888 26976 68894 26988
rect 69017 26979 69075 26985
rect 69017 26976 69029 26979
rect 68888 26948 69029 26976
rect 68888 26936 68894 26948
rect 69017 26945 69029 26948
rect 69063 26945 69075 26979
rect 69017 26939 69075 26945
rect 69106 26936 69112 26988
rect 69164 26976 69170 26988
rect 70121 26979 70179 26985
rect 69164 26948 69980 26976
rect 69164 26936 69170 26948
rect 69842 26908 69848 26920
rect 65720 26880 69848 26908
rect 65720 26849 65748 26880
rect 69842 26868 69848 26880
rect 69900 26868 69906 26920
rect 69952 26908 69980 26948
rect 70121 26945 70133 26979
rect 70167 26976 70179 26979
rect 70670 26976 70676 26988
rect 70167 26948 70676 26976
rect 70167 26945 70179 26948
rect 70121 26939 70179 26945
rect 70670 26936 70676 26948
rect 70728 26936 70734 26988
rect 70946 26976 70952 26988
rect 70907 26948 70952 26976
rect 70946 26936 70952 26948
rect 71004 26936 71010 26988
rect 72237 26979 72295 26985
rect 72237 26945 72249 26979
rect 72283 26976 72295 26979
rect 72602 26976 72608 26988
rect 72283 26948 72608 26976
rect 72283 26945 72295 26948
rect 72237 26939 72295 26945
rect 72602 26936 72608 26948
rect 72660 26936 72666 26988
rect 72329 26911 72387 26917
rect 72329 26908 72341 26911
rect 69952 26880 72341 26908
rect 72329 26877 72341 26880
rect 72375 26877 72387 26911
rect 72329 26871 72387 26877
rect 72513 26911 72571 26917
rect 72513 26877 72525 26911
rect 72559 26877 72571 26911
rect 72712 26908 72740 27016
rect 73632 27016 74580 27044
rect 73154 26976 73160 26988
rect 73115 26948 73160 26976
rect 73154 26936 73160 26948
rect 73212 26936 73218 26988
rect 73632 26985 73660 27016
rect 73617 26979 73675 26985
rect 73617 26945 73629 26979
rect 73663 26945 73675 26979
rect 73617 26939 73675 26945
rect 74261 26979 74319 26985
rect 74261 26945 74273 26979
rect 74307 26976 74319 26979
rect 74442 26976 74448 26988
rect 74307 26948 74448 26976
rect 74307 26945 74319 26948
rect 74261 26939 74319 26945
rect 74442 26936 74448 26948
rect 74500 26936 74506 26988
rect 74552 26976 74580 27016
rect 74994 27004 75000 27056
rect 75052 27044 75058 27056
rect 76009 27047 76067 27053
rect 76009 27044 76021 27047
rect 75052 27016 76021 27044
rect 75052 27004 75058 27016
rect 76009 27013 76021 27016
rect 76055 27013 76067 27047
rect 76116 27044 76144 27084
rect 77021 27081 77033 27115
rect 77067 27081 77079 27115
rect 77021 27075 77079 27081
rect 76558 27044 76564 27056
rect 76116 27016 76564 27044
rect 76009 27007 76067 27013
rect 76558 27004 76564 27016
rect 76616 27004 76622 27056
rect 77036 27044 77064 27075
rect 77294 27072 77300 27124
rect 77352 27112 77358 27124
rect 77389 27115 77447 27121
rect 77389 27112 77401 27115
rect 77352 27084 77401 27112
rect 77352 27072 77358 27084
rect 77389 27081 77401 27084
rect 77435 27081 77447 27115
rect 77389 27075 77447 27081
rect 77496 27084 78720 27112
rect 77496 27044 77524 27084
rect 77036 27016 77524 27044
rect 74552 26948 74764 26976
rect 73341 26911 73399 26917
rect 73341 26908 73353 26911
rect 72712 26880 73353 26908
rect 72513 26871 72571 26877
rect 73341 26877 73353 26880
rect 73387 26877 73399 26911
rect 74736 26908 74764 26948
rect 74810 26936 74816 26988
rect 74868 26976 74874 26988
rect 78692 26985 78720 27084
rect 79226 27072 79232 27124
rect 79284 27112 79290 27124
rect 79781 27115 79839 27121
rect 79781 27112 79793 27115
rect 79284 27084 79793 27112
rect 79284 27072 79290 27084
rect 79781 27081 79793 27084
rect 79827 27081 79839 27115
rect 79781 27075 79839 27081
rect 79870 27072 79876 27124
rect 79928 27112 79934 27124
rect 83918 27112 83924 27124
rect 79928 27084 83924 27112
rect 79928 27072 79934 27084
rect 83918 27072 83924 27084
rect 83976 27072 83982 27124
rect 84194 27072 84200 27124
rect 84252 27112 84258 27124
rect 84749 27115 84807 27121
rect 84749 27112 84761 27115
rect 84252 27084 84761 27112
rect 84252 27072 84258 27084
rect 84749 27081 84761 27084
rect 84795 27081 84807 27115
rect 84749 27075 84807 27081
rect 84930 27072 84936 27124
rect 84988 27112 84994 27124
rect 89070 27112 89076 27124
rect 84988 27084 89076 27112
rect 84988 27072 84994 27084
rect 89070 27072 89076 27084
rect 89128 27072 89134 27124
rect 90361 27115 90419 27121
rect 90361 27112 90373 27115
rect 89686 27084 90373 27112
rect 85666 27004 85672 27056
rect 85724 27044 85730 27056
rect 85724 27016 86908 27044
rect 85724 27004 85730 27016
rect 76653 26979 76711 26985
rect 77481 26980 77539 26985
rect 76653 26976 76665 26979
rect 74868 26948 76665 26976
rect 74868 26936 74874 26948
rect 76653 26945 76665 26948
rect 76699 26976 76711 26979
rect 77404 26979 77539 26980
rect 77404 26976 77493 26979
rect 76699 26952 77493 26976
rect 76699 26948 77432 26952
rect 76699 26945 76711 26948
rect 76653 26939 76711 26945
rect 77481 26945 77493 26952
rect 77527 26976 77539 26979
rect 78125 26979 78183 26985
rect 78125 26976 78137 26979
rect 77527 26948 78137 26976
rect 77527 26945 77539 26948
rect 77481 26939 77539 26945
rect 78125 26945 78137 26948
rect 78171 26945 78183 26979
rect 78125 26939 78183 26945
rect 78677 26979 78735 26985
rect 78677 26945 78689 26979
rect 78723 26945 78735 26979
rect 78677 26939 78735 26945
rect 79042 26936 79048 26988
rect 79100 26976 79106 26988
rect 79321 26979 79379 26985
rect 79321 26976 79333 26979
rect 79100 26948 79333 26976
rect 79100 26936 79106 26948
rect 79321 26945 79333 26948
rect 79367 26945 79379 26979
rect 79321 26939 79379 26945
rect 79520 26976 79732 26980
rect 79965 26979 80023 26985
rect 79965 26976 79977 26979
rect 79520 26952 79977 26976
rect 75914 26908 75920 26920
rect 74736 26880 75920 26908
rect 73341 26871 73399 26877
rect 65705 26843 65763 26849
rect 65705 26809 65717 26843
rect 65751 26809 65763 26843
rect 65705 26803 65763 26809
rect 66349 26843 66407 26849
rect 66349 26809 66361 26843
rect 66395 26840 66407 26843
rect 70302 26840 70308 26852
rect 66395 26812 70308 26840
rect 66395 26809 66407 26812
rect 66349 26803 66407 26809
rect 70302 26800 70308 26812
rect 70360 26800 70366 26852
rect 71866 26840 71872 26852
rect 71827 26812 71872 26840
rect 71866 26800 71872 26812
rect 71924 26800 71930 26852
rect 72528 26784 72556 26871
rect 75914 26868 75920 26880
rect 75972 26868 75978 26920
rect 76098 26908 76104 26920
rect 76059 26880 76104 26908
rect 76098 26868 76104 26880
rect 76156 26868 76162 26920
rect 76190 26868 76196 26920
rect 76248 26908 76254 26920
rect 77573 26911 77631 26917
rect 77573 26908 77585 26911
rect 76248 26880 77585 26908
rect 76248 26868 76254 26880
rect 77573 26877 77585 26880
rect 77619 26877 77631 26911
rect 79520 26908 79548 26952
rect 79704 26948 79977 26952
rect 79965 26945 79977 26948
rect 80011 26945 80023 26979
rect 79965 26939 80023 26945
rect 80054 26936 80060 26988
rect 80112 26976 80118 26988
rect 83844 26976 83964 26980
rect 84010 26976 84016 26988
rect 80112 26952 84016 26976
rect 80112 26948 83872 26952
rect 83936 26948 84016 26952
rect 80112 26936 80118 26948
rect 84010 26936 84016 26948
rect 84068 26985 84074 26988
rect 84068 26979 84127 26985
rect 84068 26945 84081 26979
rect 84115 26976 84127 26979
rect 84933 26979 84991 26985
rect 84115 26948 84161 26976
rect 84115 26945 84127 26948
rect 84068 26939 84127 26945
rect 84933 26945 84945 26979
rect 84979 26976 84991 26979
rect 84979 26948 85068 26976
rect 84979 26945 84991 26948
rect 84933 26939 84991 26945
rect 84068 26936 84074 26939
rect 84838 26908 84844 26920
rect 77573 26871 77631 26877
rect 79152 26880 79548 26908
rect 84166 26880 84844 26908
rect 74491 26843 74549 26849
rect 74491 26809 74503 26843
rect 74537 26840 74549 26843
rect 78674 26840 78680 26852
rect 74537 26812 78680 26840
rect 74537 26809 74549 26812
rect 74491 26803 74549 26809
rect 78674 26800 78680 26812
rect 78732 26800 78738 26852
rect 79152 26849 79180 26880
rect 79137 26843 79195 26849
rect 79137 26809 79149 26843
rect 79183 26809 79195 26843
rect 84166 26840 84194 26880
rect 84838 26868 84844 26880
rect 84896 26868 84902 26920
rect 79137 26803 79195 26809
rect 79336 26812 84194 26840
rect 84289 26843 84347 26849
rect 64555 26744 65288 26772
rect 64555 26741 64567 26744
rect 64509 26735 64567 26741
rect 66254 26732 66260 26784
rect 66312 26772 66318 26784
rect 69106 26772 69112 26784
rect 66312 26744 69112 26772
rect 66312 26732 66318 26744
rect 69106 26732 69112 26744
rect 69164 26732 69170 26784
rect 69566 26732 69572 26784
rect 69624 26772 69630 26784
rect 70394 26772 70400 26784
rect 69624 26744 70400 26772
rect 69624 26732 69630 26744
rect 70394 26732 70400 26744
rect 70452 26732 70458 26784
rect 70762 26772 70768 26784
rect 70723 26744 70768 26772
rect 70762 26732 70768 26744
rect 70820 26732 70826 26784
rect 72510 26732 72516 26784
rect 72568 26732 72574 26784
rect 72694 26732 72700 26784
rect 72752 26772 72758 26784
rect 72973 26775 73031 26781
rect 72973 26772 72985 26775
rect 72752 26744 72985 26772
rect 72752 26732 72758 26744
rect 72973 26741 72985 26744
rect 73019 26741 73031 26775
rect 72973 26735 73031 26741
rect 73062 26732 73068 26784
rect 73120 26772 73126 26784
rect 75546 26772 75552 26784
rect 73120 26744 75552 26772
rect 73120 26732 73126 26744
rect 75546 26732 75552 26744
rect 75604 26732 75610 26784
rect 75641 26775 75699 26781
rect 75641 26741 75653 26775
rect 75687 26772 75699 26775
rect 76466 26772 76472 26784
rect 75687 26744 76472 26772
rect 75687 26741 75699 26744
rect 75641 26735 75699 26741
rect 76466 26732 76472 26744
rect 76524 26732 76530 26784
rect 76558 26732 76564 26784
rect 76616 26772 76622 26784
rect 78398 26772 78404 26784
rect 76616 26744 78404 26772
rect 76616 26732 76622 26744
rect 78398 26732 78404 26744
rect 78456 26732 78462 26784
rect 78493 26775 78551 26781
rect 78493 26741 78505 26775
rect 78539 26772 78551 26775
rect 79336 26772 79364 26812
rect 84289 26809 84301 26843
rect 84335 26840 84347 26843
rect 84562 26840 84568 26852
rect 84335 26812 84568 26840
rect 84335 26809 84347 26812
rect 84289 26803 84347 26809
rect 84562 26800 84568 26812
rect 84620 26800 84626 26852
rect 78539 26744 79364 26772
rect 78539 26741 78551 26744
rect 78493 26735 78551 26741
rect 79502 26732 79508 26784
rect 79560 26772 79566 26784
rect 85040 26772 85068 26948
rect 85298 26936 85304 26988
rect 85356 26976 85362 26988
rect 86880 26985 86908 27016
rect 86954 27004 86960 27056
rect 87012 27044 87018 27056
rect 89686 27044 89714 27084
rect 90361 27081 90373 27084
rect 90407 27081 90419 27115
rect 90361 27075 90419 27081
rect 90468 27084 90680 27112
rect 87012 27016 89714 27044
rect 87012 27004 87018 27016
rect 90082 27004 90088 27056
rect 90140 27044 90146 27056
rect 90468 27044 90496 27084
rect 90140 27016 90496 27044
rect 90652 27044 90680 27084
rect 90726 27072 90732 27124
rect 90784 27112 90790 27124
rect 90784 27084 92336 27112
rect 90784 27072 90790 27084
rect 92308 27044 92336 27084
rect 92474 27072 92480 27124
rect 92532 27112 92538 27124
rect 92845 27115 92903 27121
rect 92845 27112 92857 27115
rect 92532 27084 92857 27112
rect 92532 27072 92538 27084
rect 92845 27081 92857 27084
rect 92891 27081 92903 27115
rect 94501 27115 94559 27121
rect 94501 27112 94513 27115
rect 92845 27075 92903 27081
rect 92952 27084 94513 27112
rect 92952 27044 92980 27084
rect 94501 27081 94513 27084
rect 94547 27081 94559 27115
rect 94501 27075 94559 27081
rect 95234 27072 95240 27124
rect 95292 27112 95298 27124
rect 95697 27115 95755 27121
rect 95697 27112 95709 27115
rect 95292 27084 95709 27112
rect 95292 27072 95298 27084
rect 95697 27081 95709 27084
rect 95743 27081 95755 27115
rect 95697 27075 95755 27081
rect 95786 27072 95792 27124
rect 95844 27112 95850 27124
rect 99558 27112 99564 27124
rect 95844 27084 99564 27112
rect 95844 27072 95850 27084
rect 99558 27072 99564 27084
rect 99616 27072 99622 27124
rect 100570 27112 100576 27124
rect 100531 27084 100576 27112
rect 100570 27072 100576 27084
rect 100628 27072 100634 27124
rect 104618 27072 104624 27124
rect 104676 27112 104682 27124
rect 105357 27115 105415 27121
rect 105357 27112 105369 27115
rect 104676 27084 105369 27112
rect 104676 27072 104682 27084
rect 105357 27081 105369 27084
rect 105403 27081 105415 27115
rect 110046 27112 110052 27124
rect 105357 27075 105415 27081
rect 109006 27084 110052 27112
rect 94406 27044 94412 27056
rect 90652 27016 92244 27044
rect 92308 27016 92980 27044
rect 94367 27016 94412 27044
rect 90140 27004 90146 27016
rect 85577 26979 85635 26985
rect 85577 26976 85589 26979
rect 85356 26948 85589 26976
rect 85356 26936 85362 26948
rect 85577 26945 85589 26948
rect 85623 26945 85635 26979
rect 86221 26979 86279 26985
rect 86221 26976 86233 26979
rect 85577 26939 85635 26945
rect 85684 26948 86233 26976
rect 85206 26868 85212 26920
rect 85264 26908 85270 26920
rect 85684 26908 85712 26948
rect 86221 26945 86233 26948
rect 86267 26945 86279 26979
rect 86221 26939 86279 26945
rect 86865 26979 86923 26985
rect 86865 26945 86877 26979
rect 86911 26945 86923 26979
rect 89162 26976 89168 26988
rect 86865 26939 86923 26945
rect 87248 26948 89168 26976
rect 87248 26908 87276 26948
rect 89162 26936 89168 26948
rect 89220 26936 89226 26988
rect 89622 26976 89628 26988
rect 89583 26948 89628 26976
rect 89622 26936 89628 26948
rect 89680 26936 89686 26988
rect 90174 26976 90180 26988
rect 89732 26948 90180 26976
rect 89732 26908 89760 26948
rect 90174 26936 90180 26948
rect 90232 26936 90238 26988
rect 90269 26979 90327 26985
rect 90269 26945 90281 26979
rect 90315 26976 90327 26979
rect 90358 26976 90364 26988
rect 90315 26948 90364 26976
rect 90315 26945 90327 26948
rect 90269 26939 90327 26945
rect 90358 26936 90364 26948
rect 90416 26936 90422 26988
rect 90634 26976 90640 26988
rect 90560 26948 90640 26976
rect 90560 26917 90588 26948
rect 90634 26936 90640 26948
rect 90692 26936 90698 26988
rect 91370 26976 91376 26988
rect 91331 26948 91376 26976
rect 91370 26936 91376 26948
rect 91428 26936 91434 26988
rect 92216 26976 92244 27016
rect 94406 27004 94412 27016
rect 94464 27004 94470 27056
rect 94590 27004 94596 27056
rect 94648 27044 94654 27056
rect 101674 27044 101680 27056
rect 94648 27016 101680 27044
rect 94648 27004 94654 27016
rect 101674 27004 101680 27016
rect 101732 27004 101738 27056
rect 104710 27044 104716 27056
rect 104623 27016 104716 27044
rect 104710 27004 104716 27016
rect 104768 27044 104774 27056
rect 109006 27044 109034 27084
rect 110046 27072 110052 27084
rect 110104 27072 110110 27124
rect 111518 27112 111524 27124
rect 111479 27084 111524 27112
rect 111518 27072 111524 27084
rect 111576 27072 111582 27124
rect 116305 27115 116363 27121
rect 116305 27081 116317 27115
rect 116351 27112 116363 27115
rect 117222 27112 117228 27124
rect 116351 27084 117228 27112
rect 116351 27081 116363 27084
rect 116305 27075 116363 27081
rect 117222 27072 117228 27084
rect 117280 27072 117286 27124
rect 116762 27044 116768 27056
rect 104768 27016 109034 27044
rect 116723 27016 116768 27044
rect 104768 27004 104774 27016
rect 116762 27004 116768 27016
rect 116820 27044 116826 27056
rect 117409 27047 117467 27053
rect 117409 27044 117421 27047
rect 116820 27016 117421 27044
rect 116820 27004 116826 27016
rect 117409 27013 117421 27016
rect 117455 27044 117467 27047
rect 117685 27047 117743 27053
rect 117685 27044 117697 27047
rect 117455 27016 117697 27044
rect 117455 27013 117467 27016
rect 117409 27007 117467 27013
rect 117685 27013 117697 27016
rect 117731 27013 117743 27047
rect 117685 27007 117743 27013
rect 92385 26979 92443 26985
rect 92385 26976 92397 26979
rect 92216 26948 92397 26976
rect 92385 26945 92397 26948
rect 92431 26945 92443 26979
rect 92385 26939 92443 26945
rect 93029 26979 93087 26985
rect 93029 26945 93041 26979
rect 93075 26976 93087 26979
rect 94866 26976 94872 26988
rect 93075 26948 94872 26976
rect 93075 26945 93087 26948
rect 93029 26939 93087 26945
rect 94866 26936 94872 26948
rect 94924 26936 94930 26988
rect 95234 26976 95240 26988
rect 95195 26948 95240 26976
rect 95234 26936 95240 26948
rect 95292 26936 95298 26988
rect 95878 26976 95884 26988
rect 95839 26948 95884 26976
rect 95878 26936 95884 26948
rect 95936 26936 95942 26988
rect 95970 26936 95976 26988
rect 96028 26976 96034 26988
rect 100757 26979 100815 26985
rect 96028 26948 100708 26976
rect 96028 26936 96034 26948
rect 85264 26880 85712 26908
rect 86052 26880 87276 26908
rect 87340 26880 89760 26908
rect 90545 26911 90603 26917
rect 85264 26868 85270 26880
rect 86052 26849 86080 26880
rect 86037 26843 86095 26849
rect 86037 26809 86049 26843
rect 86083 26809 86095 26843
rect 86037 26803 86095 26809
rect 86126 26800 86132 26852
rect 86184 26840 86190 26852
rect 87340 26840 87368 26880
rect 90545 26877 90557 26911
rect 90591 26877 90603 26911
rect 90545 26871 90603 26877
rect 91738 26868 91744 26920
rect 91796 26908 91802 26920
rect 100680 26908 100708 26948
rect 100757 26945 100769 26979
rect 100803 26976 100815 26979
rect 100846 26976 100852 26988
rect 100803 26948 100852 26976
rect 100803 26945 100815 26948
rect 100757 26939 100815 26945
rect 100846 26936 100852 26948
rect 100904 26936 100910 26988
rect 103330 26936 103336 26988
rect 103388 26976 103394 26988
rect 103701 26979 103759 26985
rect 103701 26976 103713 26979
rect 103388 26948 103713 26976
rect 103388 26936 103394 26948
rect 103701 26945 103713 26948
rect 103747 26945 103759 26979
rect 105538 26976 105544 26988
rect 105499 26948 105544 26976
rect 103701 26939 103759 26945
rect 105538 26936 105544 26948
rect 105596 26936 105602 26988
rect 111702 26976 111708 26988
rect 111663 26948 111708 26976
rect 111702 26936 111708 26948
rect 111760 26936 111766 26988
rect 116489 26979 116547 26985
rect 116489 26945 116501 26979
rect 116535 26945 116547 26979
rect 116489 26939 116547 26945
rect 104342 26908 104348 26920
rect 91796 26880 100616 26908
rect 100680 26880 104348 26908
rect 91796 26868 91802 26880
rect 86184 26812 87368 26840
rect 89901 26843 89959 26849
rect 86184 26800 86190 26812
rect 89901 26809 89913 26843
rect 89947 26840 89959 26843
rect 91830 26840 91836 26852
rect 89947 26812 91836 26840
rect 89947 26809 89959 26812
rect 89901 26803 89959 26809
rect 91830 26800 91836 26812
rect 91888 26800 91894 26852
rect 92198 26840 92204 26852
rect 92159 26812 92204 26840
rect 92198 26800 92204 26812
rect 92256 26800 92262 26852
rect 94038 26800 94044 26852
rect 94096 26840 94102 26852
rect 95053 26843 95111 26849
rect 95053 26840 95065 26843
rect 94096 26812 95065 26840
rect 94096 26800 94102 26812
rect 95053 26809 95065 26812
rect 95099 26809 95111 26843
rect 100202 26840 100208 26852
rect 95053 26803 95111 26809
rect 95160 26812 100208 26840
rect 85390 26772 85396 26784
rect 79560 26744 85068 26772
rect 85351 26744 85396 26772
rect 79560 26732 79566 26744
rect 85390 26732 85396 26744
rect 85448 26732 85454 26784
rect 86218 26732 86224 26784
rect 86276 26772 86282 26784
rect 86681 26775 86739 26781
rect 86681 26772 86693 26775
rect 86276 26744 86693 26772
rect 86276 26732 86282 26744
rect 86681 26741 86693 26744
rect 86727 26741 86739 26775
rect 86681 26735 86739 26741
rect 86862 26732 86868 26784
rect 86920 26772 86926 26784
rect 89441 26775 89499 26781
rect 89441 26772 89453 26775
rect 86920 26744 89453 26772
rect 86920 26732 86926 26744
rect 89441 26741 89453 26744
rect 89487 26741 89499 26775
rect 89441 26735 89499 26741
rect 90082 26732 90088 26784
rect 90140 26772 90146 26784
rect 90726 26772 90732 26784
rect 90140 26744 90732 26772
rect 90140 26732 90146 26744
rect 90726 26732 90732 26744
rect 90784 26732 90790 26784
rect 90910 26772 90916 26784
rect 90871 26744 90916 26772
rect 90910 26732 90916 26744
rect 90968 26772 90974 26784
rect 91465 26775 91523 26781
rect 91465 26772 91477 26775
rect 90968 26744 91477 26772
rect 90968 26732 90974 26744
rect 91465 26741 91477 26744
rect 91511 26741 91523 26775
rect 91465 26735 91523 26741
rect 91738 26732 91744 26784
rect 91796 26772 91802 26784
rect 95160 26772 95188 26812
rect 100202 26800 100208 26812
rect 100260 26800 100266 26852
rect 100588 26840 100616 26880
rect 104342 26868 104348 26880
rect 104400 26868 104406 26920
rect 108482 26908 108488 26920
rect 104452 26880 108488 26908
rect 104452 26840 104480 26880
rect 108482 26868 108488 26880
rect 108540 26868 108546 26920
rect 109586 26868 109592 26920
rect 109644 26908 109650 26920
rect 113634 26908 113640 26920
rect 109644 26880 113640 26908
rect 109644 26868 109650 26880
rect 113634 26868 113640 26880
rect 113692 26868 113698 26920
rect 104894 26840 104900 26852
rect 100588 26812 104480 26840
rect 104855 26812 104900 26840
rect 104894 26800 104900 26812
rect 104952 26800 104958 26852
rect 116504 26840 116532 26939
rect 117130 26936 117136 26988
rect 117188 26976 117194 26988
rect 117225 26979 117283 26985
rect 117225 26976 117237 26979
rect 117188 26948 117237 26976
rect 117188 26936 117194 26948
rect 117225 26945 117237 26948
rect 117271 26945 117283 26979
rect 117958 26976 117964 26988
rect 117919 26948 117964 26976
rect 117225 26939 117283 26945
rect 117958 26936 117964 26948
rect 118016 26936 118022 26988
rect 105280 26812 116532 26840
rect 91796 26744 95188 26772
rect 103517 26775 103575 26781
rect 91796 26732 91802 26744
rect 103517 26741 103529 26775
rect 103563 26772 103575 26775
rect 105280 26772 105308 26812
rect 103563 26744 105308 26772
rect 103563 26741 103575 26744
rect 103517 26735 103575 26741
rect 117774 26732 117780 26784
rect 117832 26772 117838 26784
rect 118053 26775 118111 26781
rect 118053 26772 118065 26775
rect 117832 26744 118065 26772
rect 117832 26732 117838 26744
rect 118053 26741 118065 26744
rect 118099 26741 118111 26775
rect 118053 26735 118111 26741
rect 1104 26682 118864 26704
rect 1104 26630 15674 26682
rect 15726 26630 15738 26682
rect 15790 26630 15802 26682
rect 15854 26630 15866 26682
rect 15918 26630 15930 26682
rect 15982 26630 45122 26682
rect 45174 26630 45186 26682
rect 45238 26630 45250 26682
rect 45302 26630 45314 26682
rect 45366 26630 45378 26682
rect 45430 26630 74570 26682
rect 74622 26630 74634 26682
rect 74686 26630 74698 26682
rect 74750 26630 74762 26682
rect 74814 26630 74826 26682
rect 74878 26630 104018 26682
rect 104070 26630 104082 26682
rect 104134 26630 104146 26682
rect 104198 26630 104210 26682
rect 104262 26630 104274 26682
rect 104326 26630 118864 26682
rect 1104 26608 118864 26630
rect 1670 26528 1676 26580
rect 1728 26568 1734 26580
rect 22094 26568 22100 26580
rect 1728 26540 22100 26568
rect 1728 26528 1734 26540
rect 22094 26528 22100 26540
rect 22152 26528 22158 26580
rect 24118 26528 24124 26580
rect 24176 26568 24182 26580
rect 29546 26568 29552 26580
rect 24176 26540 29552 26568
rect 24176 26528 24182 26540
rect 29546 26528 29552 26540
rect 29604 26528 29610 26580
rect 29730 26568 29736 26580
rect 29691 26540 29736 26568
rect 29730 26528 29736 26540
rect 29788 26528 29794 26580
rect 31478 26528 31484 26580
rect 31536 26568 31542 26580
rect 40954 26568 40960 26580
rect 31536 26540 40960 26568
rect 31536 26528 31542 26540
rect 40954 26528 40960 26540
rect 41012 26528 41018 26580
rect 41230 26528 41236 26580
rect 41288 26568 41294 26580
rect 46198 26568 46204 26580
rect 41288 26540 46204 26568
rect 41288 26528 41294 26540
rect 46198 26528 46204 26540
rect 46256 26528 46262 26580
rect 46477 26571 46535 26577
rect 46477 26537 46489 26571
rect 46523 26568 46535 26571
rect 46566 26568 46572 26580
rect 46523 26540 46572 26568
rect 46523 26537 46535 26540
rect 46477 26531 46535 26537
rect 46566 26528 46572 26540
rect 46624 26528 46630 26580
rect 46750 26528 46756 26580
rect 46808 26568 46814 26580
rect 50890 26568 50896 26580
rect 46808 26540 50896 26568
rect 46808 26528 46814 26540
rect 50890 26528 50896 26540
rect 50948 26528 50954 26580
rect 51166 26528 51172 26580
rect 51224 26568 51230 26580
rect 60550 26568 60556 26580
rect 51224 26540 60556 26568
rect 51224 26528 51230 26540
rect 60550 26528 60556 26540
rect 60608 26528 60614 26580
rect 61746 26528 61752 26580
rect 61804 26568 61810 26580
rect 68370 26568 68376 26580
rect 61804 26540 68376 26568
rect 61804 26528 61810 26540
rect 68370 26528 68376 26540
rect 68428 26528 68434 26580
rect 68462 26528 68468 26580
rect 68520 26568 68526 26580
rect 69109 26571 69167 26577
rect 69109 26568 69121 26571
rect 68520 26540 69121 26568
rect 68520 26528 68526 26540
rect 69109 26537 69121 26540
rect 69155 26537 69167 26571
rect 70026 26568 70032 26580
rect 69987 26540 70032 26568
rect 69109 26531 69167 26537
rect 70026 26528 70032 26540
rect 70084 26528 70090 26580
rect 70366 26540 74856 26568
rect 2685 26503 2743 26509
rect 2685 26469 2697 26503
rect 2731 26500 2743 26503
rect 2774 26500 2780 26512
rect 2731 26472 2780 26500
rect 2731 26469 2743 26472
rect 2685 26463 2743 26469
rect 2774 26460 2780 26472
rect 2832 26460 2838 26512
rect 15562 26460 15568 26512
rect 15620 26500 15626 26512
rect 21174 26500 21180 26512
rect 15620 26472 21180 26500
rect 15620 26460 15626 26472
rect 21174 26460 21180 26472
rect 21232 26460 21238 26512
rect 22370 26460 22376 26512
rect 22428 26500 22434 26512
rect 30098 26500 30104 26512
rect 22428 26472 30104 26500
rect 22428 26460 22434 26472
rect 30098 26460 30104 26472
rect 30156 26460 30162 26512
rect 30190 26460 30196 26512
rect 30248 26500 30254 26512
rect 31754 26500 31760 26512
rect 30248 26472 31760 26500
rect 30248 26460 30254 26472
rect 31754 26460 31760 26472
rect 31812 26460 31818 26512
rect 31846 26460 31852 26512
rect 31904 26500 31910 26512
rect 43438 26500 43444 26512
rect 31904 26472 43444 26500
rect 31904 26460 31910 26472
rect 43438 26460 43444 26472
rect 43496 26460 43502 26512
rect 45646 26460 45652 26512
rect 45704 26500 45710 26512
rect 48222 26500 48228 26512
rect 45704 26472 48228 26500
rect 45704 26460 45710 26472
rect 48222 26460 48228 26472
rect 48280 26460 48286 26512
rect 49053 26503 49111 26509
rect 49053 26469 49065 26503
rect 49099 26500 49111 26503
rect 50798 26500 50804 26512
rect 49099 26472 50804 26500
rect 49099 26469 49111 26472
rect 49053 26463 49111 26469
rect 50798 26460 50804 26472
rect 50856 26460 50862 26512
rect 50908 26472 51074 26500
rect 1210 26392 1216 26444
rect 1268 26432 1274 26444
rect 1397 26435 1455 26441
rect 1397 26432 1409 26435
rect 1268 26404 1409 26432
rect 1268 26392 1274 26404
rect 1397 26401 1409 26404
rect 1443 26401 1455 26435
rect 1397 26395 1455 26401
rect 6638 26392 6644 26444
rect 6696 26432 6702 26444
rect 24118 26432 24124 26444
rect 6696 26404 24124 26432
rect 6696 26392 6702 26404
rect 24118 26392 24124 26404
rect 24176 26392 24182 26444
rect 28166 26392 28172 26444
rect 28224 26432 28230 26444
rect 31570 26432 31576 26444
rect 28224 26404 31576 26432
rect 28224 26392 28230 26404
rect 31570 26392 31576 26404
rect 31628 26392 31634 26444
rect 31662 26392 31668 26444
rect 31720 26432 31726 26444
rect 35802 26432 35808 26444
rect 31720 26404 35664 26432
rect 35763 26404 35808 26432
rect 31720 26392 31726 26404
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26333 1731 26367
rect 1673 26327 1731 26333
rect 2869 26367 2927 26373
rect 2869 26333 2881 26367
rect 2915 26364 2927 26367
rect 22370 26364 22376 26376
rect 2915 26336 22376 26364
rect 2915 26333 2927 26336
rect 2869 26327 2927 26333
rect 1688 26296 1716 26327
rect 22370 26324 22376 26336
rect 22428 26324 22434 26376
rect 29454 26364 29460 26376
rect 24412 26336 29460 26364
rect 1688 26268 19334 26296
rect 14 26188 20 26240
rect 72 26228 78 26240
rect 2866 26228 2872 26240
rect 72 26200 2872 26228
rect 72 26188 78 26200
rect 2866 26188 2872 26200
rect 2924 26188 2930 26240
rect 9030 26188 9036 26240
rect 9088 26228 9094 26240
rect 10318 26228 10324 26240
rect 9088 26200 10324 26228
rect 9088 26188 9094 26200
rect 10318 26188 10324 26200
rect 10376 26188 10382 26240
rect 19306 26228 19334 26268
rect 24412 26228 24440 26336
rect 29454 26324 29460 26336
rect 29512 26324 29518 26376
rect 29638 26324 29644 26376
rect 29696 26364 29702 26376
rect 29917 26367 29975 26373
rect 29917 26364 29929 26367
rect 29696 26336 29929 26364
rect 29696 26324 29702 26336
rect 29917 26333 29929 26336
rect 29963 26333 29975 26367
rect 35526 26364 35532 26376
rect 29917 26327 29975 26333
rect 30024 26336 35532 26364
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 30024 26296 30052 26336
rect 35526 26324 35532 26336
rect 35584 26324 35590 26376
rect 35636 26364 35664 26404
rect 35802 26392 35808 26404
rect 35860 26392 35866 26444
rect 35894 26392 35900 26444
rect 35952 26432 35958 26444
rect 40770 26432 40776 26444
rect 35952 26404 40776 26432
rect 35952 26392 35958 26404
rect 40770 26392 40776 26404
rect 40828 26392 40834 26444
rect 41230 26392 41236 26444
rect 41288 26432 41294 26444
rect 50908 26432 50936 26472
rect 41288 26404 41460 26432
rect 41288 26392 41294 26404
rect 41046 26364 41052 26376
rect 35636 26336 41052 26364
rect 41046 26324 41052 26336
rect 41104 26324 41110 26376
rect 41432 26364 41460 26404
rect 41616 26404 50936 26432
rect 51046 26432 51074 26472
rect 51442 26460 51448 26512
rect 51500 26500 51506 26512
rect 53561 26503 53619 26509
rect 53561 26500 53573 26503
rect 51500 26472 53573 26500
rect 51500 26460 51506 26472
rect 53561 26469 53573 26472
rect 53607 26469 53619 26503
rect 53561 26463 53619 26469
rect 54573 26503 54631 26509
rect 54573 26469 54585 26503
rect 54619 26500 54631 26503
rect 54754 26500 54760 26512
rect 54619 26472 54760 26500
rect 54619 26469 54631 26472
rect 54573 26463 54631 26469
rect 54754 26460 54760 26472
rect 54812 26460 54818 26512
rect 55309 26503 55367 26509
rect 55309 26469 55321 26503
rect 55355 26500 55367 26503
rect 56318 26500 56324 26512
rect 55355 26472 56324 26500
rect 55355 26469 55367 26472
rect 55309 26463 55367 26469
rect 56318 26460 56324 26472
rect 56376 26460 56382 26512
rect 56413 26503 56471 26509
rect 56413 26469 56425 26503
rect 56459 26500 56471 26503
rect 57330 26500 57336 26512
rect 56459 26472 57336 26500
rect 56459 26469 56471 26472
rect 56413 26463 56471 26469
rect 57330 26460 57336 26472
rect 57388 26460 57394 26512
rect 58710 26500 58716 26512
rect 58671 26472 58716 26500
rect 58710 26460 58716 26472
rect 58768 26460 58774 26512
rect 70366 26500 70394 26540
rect 61672 26472 70394 26500
rect 54386 26432 54392 26444
rect 51046 26404 54392 26432
rect 41616 26364 41644 26404
rect 54386 26392 54392 26404
rect 54444 26392 54450 26444
rect 61672 26432 61700 26472
rect 70486 26460 70492 26512
rect 70544 26500 70550 26512
rect 74718 26500 74724 26512
rect 70544 26472 74724 26500
rect 70544 26460 70550 26472
rect 74718 26460 74724 26472
rect 74776 26460 74782 26512
rect 74828 26500 74856 26540
rect 74902 26528 74908 26580
rect 74960 26568 74966 26580
rect 76558 26568 76564 26580
rect 74960 26540 76564 26568
rect 74960 26528 74966 26540
rect 76558 26528 76564 26540
rect 76616 26528 76622 26580
rect 77386 26568 77392 26580
rect 77347 26540 77392 26568
rect 77386 26528 77392 26540
rect 77444 26528 77450 26580
rect 78398 26528 78404 26580
rect 78456 26568 78462 26580
rect 79502 26568 79508 26580
rect 78456 26540 79508 26568
rect 78456 26528 78462 26540
rect 79502 26528 79508 26540
rect 79560 26528 79566 26580
rect 79612 26540 81112 26568
rect 74828 26472 77616 26500
rect 54772 26404 61700 26432
rect 46658 26364 46664 26376
rect 41432 26336 41644 26364
rect 46619 26336 46664 26364
rect 46658 26324 46664 26336
rect 46716 26324 46722 26376
rect 48222 26364 48228 26376
rect 48183 26336 48228 26364
rect 48222 26324 48228 26336
rect 48280 26324 48286 26376
rect 49234 26364 49240 26376
rect 49195 26336 49240 26364
rect 49234 26324 49240 26336
rect 49292 26324 49298 26376
rect 50338 26324 50344 26376
rect 50396 26364 50402 26376
rect 53742 26364 53748 26376
rect 50396 26336 50441 26364
rect 53703 26336 53748 26364
rect 50396 26324 50402 26336
rect 53742 26324 53748 26336
rect 53800 26324 53806 26376
rect 54772 26373 54800 26404
rect 61746 26392 61752 26444
rect 61804 26432 61810 26444
rect 61841 26435 61899 26441
rect 61841 26432 61853 26435
rect 61804 26404 61853 26432
rect 61804 26392 61810 26404
rect 61841 26401 61853 26404
rect 61887 26401 61899 26435
rect 61841 26395 61899 26401
rect 61948 26404 62804 26432
rect 54757 26367 54815 26373
rect 54757 26333 54769 26367
rect 54803 26333 54815 26367
rect 54757 26327 54815 26333
rect 55493 26367 55551 26373
rect 55493 26333 55505 26367
rect 55539 26364 55551 26367
rect 56597 26367 56655 26373
rect 56597 26364 56609 26367
rect 55539 26336 56609 26364
rect 55539 26333 55551 26336
rect 55493 26327 55551 26333
rect 56597 26333 56609 26336
rect 56643 26333 56655 26367
rect 56597 26327 56655 26333
rect 24544 26268 30052 26296
rect 24544 26256 24550 26268
rect 30098 26256 30104 26308
rect 30156 26296 30162 26308
rect 31754 26296 31760 26308
rect 30156 26268 31760 26296
rect 30156 26256 30162 26268
rect 31754 26256 31760 26268
rect 31812 26256 31818 26308
rect 35621 26299 35679 26305
rect 35621 26296 35633 26299
rect 31864 26268 35633 26296
rect 19306 26200 24440 26228
rect 26786 26188 26792 26240
rect 26844 26228 26850 26240
rect 31864 26228 31892 26268
rect 35621 26265 35633 26268
rect 35667 26265 35679 26299
rect 35621 26259 35679 26265
rect 35710 26256 35716 26308
rect 35768 26296 35774 26308
rect 40954 26296 40960 26308
rect 35768 26268 40960 26296
rect 35768 26256 35774 26268
rect 40954 26256 40960 26268
rect 41012 26256 41018 26308
rect 41414 26256 41420 26308
rect 41472 26296 41478 26308
rect 46842 26296 46848 26308
rect 41472 26268 46848 26296
rect 41472 26256 41478 26268
rect 46842 26256 46848 26268
rect 46900 26256 46906 26308
rect 47302 26256 47308 26308
rect 47360 26296 47366 26308
rect 50982 26296 50988 26308
rect 47360 26268 50988 26296
rect 47360 26256 47366 26268
rect 50982 26256 50988 26268
rect 51040 26256 51046 26308
rect 51258 26256 51264 26308
rect 51316 26296 51322 26308
rect 53374 26296 53380 26308
rect 51316 26268 53380 26296
rect 51316 26256 51322 26268
rect 53374 26256 53380 26268
rect 53432 26256 53438 26308
rect 53558 26256 53564 26308
rect 53616 26296 53622 26308
rect 55508 26296 55536 26327
rect 56870 26324 56876 26376
rect 56928 26364 56934 26376
rect 58897 26367 58955 26373
rect 58897 26364 58909 26367
rect 56928 26336 58909 26364
rect 56928 26324 56934 26336
rect 58897 26333 58909 26336
rect 58943 26333 58955 26367
rect 61010 26364 61016 26376
rect 58897 26327 58955 26333
rect 59096 26336 61016 26364
rect 59096 26296 59124 26336
rect 61010 26324 61016 26336
rect 61068 26324 61074 26376
rect 61102 26324 61108 26376
rect 61160 26364 61166 26376
rect 61948 26364 61976 26404
rect 62669 26367 62727 26373
rect 62669 26364 62681 26367
rect 61160 26336 61976 26364
rect 62040 26336 62681 26364
rect 61160 26324 61166 26336
rect 53616 26268 55536 26296
rect 55600 26268 59124 26296
rect 53616 26256 53622 26268
rect 35158 26228 35164 26240
rect 26844 26200 31892 26228
rect 35119 26200 35164 26228
rect 26844 26188 26850 26200
rect 35158 26188 35164 26200
rect 35216 26188 35222 26240
rect 35342 26188 35348 26240
rect 35400 26228 35406 26240
rect 35529 26231 35587 26237
rect 35529 26228 35541 26231
rect 35400 26200 35541 26228
rect 35400 26188 35406 26200
rect 35529 26197 35541 26200
rect 35575 26197 35587 26231
rect 35529 26191 35587 26197
rect 37642 26188 37648 26240
rect 37700 26228 37706 26240
rect 40218 26228 40224 26240
rect 37700 26200 40224 26228
rect 37700 26188 37706 26200
rect 40218 26188 40224 26200
rect 40276 26188 40282 26240
rect 48041 26231 48099 26237
rect 48041 26197 48053 26231
rect 48087 26228 48099 26231
rect 49970 26228 49976 26240
rect 48087 26200 49976 26228
rect 48087 26197 48099 26200
rect 48041 26191 48099 26197
rect 49970 26188 49976 26200
rect 50028 26188 50034 26240
rect 50154 26228 50160 26240
rect 50115 26200 50160 26228
rect 50154 26188 50160 26200
rect 50212 26188 50218 26240
rect 50522 26188 50528 26240
rect 50580 26228 50586 26240
rect 55600 26228 55628 26268
rect 59170 26256 59176 26308
rect 59228 26296 59234 26308
rect 60734 26296 60740 26308
rect 59228 26268 60740 26296
rect 59228 26256 59234 26268
rect 60734 26256 60740 26268
rect 60792 26256 60798 26308
rect 61657 26299 61715 26305
rect 61657 26296 61669 26299
rect 60844 26268 61669 26296
rect 50580 26200 55628 26228
rect 50580 26188 50586 26200
rect 55674 26188 55680 26240
rect 55732 26228 55738 26240
rect 60458 26228 60464 26240
rect 55732 26200 60464 26228
rect 55732 26188 55738 26200
rect 60458 26188 60464 26200
rect 60516 26188 60522 26240
rect 60550 26188 60556 26240
rect 60608 26228 60614 26240
rect 60844 26228 60872 26268
rect 61657 26265 61669 26268
rect 61703 26265 61715 26299
rect 61657 26259 61715 26265
rect 61749 26299 61807 26305
rect 61749 26265 61761 26299
rect 61795 26296 61807 26299
rect 61930 26296 61936 26308
rect 61795 26268 61936 26296
rect 61795 26265 61807 26268
rect 61749 26259 61807 26265
rect 61930 26256 61936 26268
rect 61988 26256 61994 26308
rect 60608 26200 60872 26228
rect 61289 26231 61347 26237
rect 60608 26188 60614 26200
rect 61289 26197 61301 26231
rect 61335 26228 61347 26231
rect 62040 26228 62068 26336
rect 62669 26333 62681 26336
rect 62715 26333 62727 26367
rect 62776 26364 62804 26404
rect 63494 26392 63500 26444
rect 63552 26432 63558 26444
rect 69934 26432 69940 26444
rect 63552 26404 69940 26432
rect 63552 26392 63558 26404
rect 69934 26392 69940 26404
rect 69992 26392 69998 26444
rect 70872 26404 72188 26432
rect 68554 26364 68560 26376
rect 62776 26336 68560 26364
rect 62669 26327 62727 26333
rect 68554 26324 68560 26336
rect 68612 26324 68618 26376
rect 68646 26324 68652 26376
rect 68704 26364 68710 26376
rect 69293 26367 69351 26373
rect 69293 26364 69305 26367
rect 68704 26336 69305 26364
rect 68704 26324 68710 26336
rect 69293 26333 69305 26336
rect 69339 26333 69351 26367
rect 69293 26327 69351 26333
rect 70213 26367 70271 26373
rect 70213 26333 70225 26367
rect 70259 26364 70271 26367
rect 70762 26364 70768 26376
rect 70259 26360 70440 26364
rect 70504 26360 70768 26364
rect 70259 26336 70768 26360
rect 70259 26333 70271 26336
rect 70213 26327 70271 26333
rect 70412 26332 70532 26336
rect 70762 26324 70768 26336
rect 70820 26324 70826 26376
rect 70872 26296 70900 26404
rect 71774 26324 71780 26376
rect 71832 26364 71838 26376
rect 72053 26367 72111 26373
rect 72053 26364 72065 26367
rect 71832 26336 72065 26364
rect 71832 26324 71838 26336
rect 72053 26333 72065 26336
rect 72099 26333 72111 26367
rect 72160 26364 72188 26404
rect 72234 26392 72240 26444
rect 72292 26432 72298 26444
rect 77478 26432 77484 26444
rect 72292 26404 77484 26432
rect 72292 26392 72298 26404
rect 77478 26392 77484 26404
rect 77536 26392 77542 26444
rect 77588 26432 77616 26472
rect 79042 26460 79048 26512
rect 79100 26500 79106 26512
rect 79137 26503 79195 26509
rect 79137 26500 79149 26503
rect 79100 26472 79149 26500
rect 79100 26460 79106 26472
rect 79137 26469 79149 26472
rect 79183 26469 79195 26503
rect 79137 26463 79195 26469
rect 79612 26432 79640 26540
rect 81084 26500 81112 26540
rect 84010 26528 84016 26580
rect 84068 26568 84074 26580
rect 85298 26568 85304 26580
rect 84068 26540 85304 26568
rect 84068 26528 84074 26540
rect 85298 26528 85304 26540
rect 85356 26528 85362 26580
rect 85390 26528 85396 26580
rect 85448 26568 85454 26580
rect 100846 26568 100852 26580
rect 85448 26540 100852 26568
rect 85448 26528 85454 26540
rect 100846 26528 100852 26540
rect 100904 26528 100910 26580
rect 104342 26528 104348 26580
rect 104400 26568 104406 26580
rect 110966 26568 110972 26580
rect 104400 26540 110972 26568
rect 104400 26528 104406 26540
rect 110966 26528 110972 26540
rect 111024 26528 111030 26580
rect 90082 26500 90088 26512
rect 81084 26472 90088 26500
rect 90082 26460 90088 26472
rect 90140 26460 90146 26512
rect 90284 26472 95740 26500
rect 77588 26404 79640 26432
rect 79781 26435 79839 26441
rect 79781 26401 79793 26435
rect 79827 26401 79839 26435
rect 79781 26395 79839 26401
rect 74902 26364 74908 26376
rect 72160 26336 74908 26364
rect 72053 26327 72111 26333
rect 74902 26324 74908 26336
rect 74960 26324 74966 26376
rect 74997 26367 75055 26373
rect 74997 26333 75009 26367
rect 75043 26364 75055 26367
rect 75086 26364 75092 26376
rect 75043 26336 75092 26364
rect 75043 26333 75055 26336
rect 74997 26327 75055 26333
rect 75086 26324 75092 26336
rect 75144 26324 75150 26376
rect 76466 26364 76472 26376
rect 76427 26336 76472 26364
rect 76466 26324 76472 26336
rect 76524 26324 76530 26376
rect 77570 26364 77576 26376
rect 77531 26336 77576 26364
rect 77570 26324 77576 26336
rect 77628 26324 77634 26376
rect 78674 26324 78680 26376
rect 78732 26364 78738 26376
rect 78732 26336 79640 26364
rect 78732 26324 78738 26336
rect 71225 26299 71283 26305
rect 71225 26296 71237 26299
rect 62500 26268 70900 26296
rect 70964 26268 71237 26296
rect 62500 26237 62528 26268
rect 61335 26200 62068 26228
rect 62485 26231 62543 26237
rect 61335 26197 61347 26200
rect 61289 26191 61347 26197
rect 62485 26197 62497 26231
rect 62531 26197 62543 26231
rect 62485 26191 62543 26197
rect 70670 26188 70676 26240
rect 70728 26228 70734 26240
rect 70964 26228 70992 26268
rect 71225 26265 71237 26268
rect 71271 26296 71283 26299
rect 71314 26296 71320 26308
rect 71271 26268 71320 26296
rect 71271 26265 71283 26268
rect 71225 26259 71283 26265
rect 71314 26256 71320 26268
rect 71372 26256 71378 26308
rect 71409 26299 71467 26305
rect 71409 26265 71421 26299
rect 71455 26296 71467 26299
rect 71590 26296 71596 26308
rect 71455 26268 71596 26296
rect 71455 26265 71467 26268
rect 71409 26259 71467 26265
rect 71590 26256 71596 26268
rect 71648 26256 71654 26308
rect 72786 26256 72792 26308
rect 72844 26296 72850 26308
rect 79505 26299 79563 26305
rect 79505 26296 79517 26299
rect 72844 26268 79517 26296
rect 72844 26256 72850 26268
rect 79505 26265 79517 26268
rect 79551 26265 79563 26299
rect 79612 26296 79640 26336
rect 79686 26324 79692 26376
rect 79744 26364 79750 26376
rect 79796 26364 79824 26395
rect 82262 26392 82268 26444
rect 82320 26432 82326 26444
rect 82320 26404 90128 26432
rect 82320 26392 82326 26404
rect 79744 26336 79824 26364
rect 79744 26324 79750 26336
rect 81894 26324 81900 26376
rect 81952 26364 81958 26376
rect 89070 26364 89076 26376
rect 81952 26336 89076 26364
rect 81952 26324 81958 26336
rect 89070 26324 89076 26336
rect 89128 26324 89134 26376
rect 89990 26364 89996 26376
rect 89272 26336 89996 26364
rect 79612 26268 79732 26296
rect 79505 26259 79563 26265
rect 70728 26200 70992 26228
rect 70728 26188 70734 26200
rect 71038 26188 71044 26240
rect 71096 26228 71102 26240
rect 71774 26228 71780 26240
rect 71096 26200 71780 26228
rect 71096 26188 71102 26200
rect 71774 26188 71780 26200
rect 71832 26188 71838 26240
rect 71866 26188 71872 26240
rect 71924 26228 71930 26240
rect 71924 26200 71969 26228
rect 71924 26188 71930 26200
rect 74718 26188 74724 26240
rect 74776 26228 74782 26240
rect 74813 26231 74871 26237
rect 74813 26228 74825 26231
rect 74776 26200 74825 26228
rect 74776 26188 74782 26200
rect 74813 26197 74825 26200
rect 74859 26197 74871 26231
rect 76650 26228 76656 26240
rect 76611 26200 76656 26228
rect 74813 26191 74871 26197
rect 76650 26188 76656 26200
rect 76708 26188 76714 26240
rect 79594 26228 79600 26240
rect 79555 26200 79600 26228
rect 79594 26188 79600 26200
rect 79652 26188 79658 26240
rect 79704 26228 79732 26268
rect 81158 26256 81164 26308
rect 81216 26296 81222 26308
rect 89162 26296 89168 26308
rect 81216 26268 89168 26296
rect 81216 26256 81222 26268
rect 89162 26256 89168 26268
rect 89220 26256 89226 26308
rect 89272 26228 89300 26336
rect 89990 26324 89996 26336
rect 90048 26324 90054 26376
rect 90100 26364 90128 26404
rect 90174 26392 90180 26444
rect 90232 26432 90238 26444
rect 90284 26432 90312 26472
rect 91738 26432 91744 26444
rect 90232 26404 90312 26432
rect 90376 26404 91744 26432
rect 90232 26392 90238 26404
rect 90376 26364 90404 26404
rect 91738 26392 91744 26404
rect 91796 26392 91802 26444
rect 92017 26435 92075 26441
rect 92017 26401 92029 26435
rect 92063 26432 92075 26435
rect 95712 26432 95740 26472
rect 95786 26460 95792 26512
rect 95844 26500 95850 26512
rect 103330 26500 103336 26512
rect 95844 26472 103336 26500
rect 95844 26460 95850 26472
rect 103330 26460 103336 26472
rect 103388 26460 103394 26512
rect 117317 26503 117375 26509
rect 117317 26469 117329 26503
rect 117363 26500 117375 26503
rect 117406 26500 117412 26512
rect 117363 26472 117412 26500
rect 117363 26469 117375 26472
rect 117317 26463 117375 26469
rect 117406 26460 117412 26472
rect 117464 26460 117470 26512
rect 102778 26432 102784 26444
rect 92063 26404 95648 26432
rect 95712 26404 102784 26432
rect 92063 26401 92075 26404
rect 92017 26395 92075 26401
rect 90100 26336 90404 26364
rect 90450 26324 90456 26376
rect 90508 26364 90514 26376
rect 93670 26364 93676 26376
rect 90508 26336 90553 26364
rect 90652 26336 92244 26364
rect 93631 26336 93676 26364
rect 90508 26324 90514 26336
rect 89346 26256 89352 26308
rect 89404 26296 89410 26308
rect 89404 26268 90404 26296
rect 89404 26256 89410 26268
rect 90266 26228 90272 26240
rect 79704 26200 89300 26228
rect 90227 26200 90272 26228
rect 90266 26188 90272 26200
rect 90324 26188 90330 26240
rect 90376 26228 90404 26268
rect 90652 26228 90680 26336
rect 91830 26256 91836 26308
rect 91888 26296 91894 26308
rect 92216 26296 92244 26336
rect 93670 26324 93676 26336
rect 93728 26324 93734 26376
rect 95620 26364 95648 26404
rect 102778 26392 102784 26404
rect 102836 26392 102842 26444
rect 116854 26364 116860 26376
rect 95620 26336 116860 26364
rect 116854 26324 116860 26336
rect 116912 26324 116918 26376
rect 117038 26324 117044 26376
rect 117096 26364 117102 26376
rect 117133 26367 117191 26373
rect 117133 26364 117145 26367
rect 117096 26336 117145 26364
rect 117096 26324 117102 26336
rect 117133 26333 117145 26336
rect 117179 26333 117191 26367
rect 117133 26327 117191 26333
rect 117961 26367 118019 26373
rect 117961 26333 117973 26367
rect 118007 26364 118019 26367
rect 118510 26364 118516 26376
rect 118007 26336 118516 26364
rect 118007 26333 118019 26336
rect 117961 26327 118019 26333
rect 118510 26324 118516 26336
rect 118568 26324 118574 26376
rect 117774 26296 117780 26308
rect 91888 26268 91933 26296
rect 92216 26268 117780 26296
rect 91888 26256 91894 26268
rect 117774 26256 117780 26268
rect 117832 26256 117838 26308
rect 118050 26256 118056 26308
rect 118108 26296 118114 26308
rect 118145 26299 118203 26305
rect 118145 26296 118157 26299
rect 118108 26268 118157 26296
rect 118108 26256 118114 26268
rect 118145 26265 118157 26268
rect 118191 26265 118203 26299
rect 118145 26259 118203 26265
rect 93486 26228 93492 26240
rect 90376 26200 90680 26228
rect 93447 26200 93492 26228
rect 93486 26188 93492 26200
rect 93544 26188 93550 26240
rect 1104 26138 118864 26160
rect 1104 26086 30398 26138
rect 30450 26086 30462 26138
rect 30514 26086 30526 26138
rect 30578 26086 30590 26138
rect 30642 26086 30654 26138
rect 30706 26086 59846 26138
rect 59898 26086 59910 26138
rect 59962 26086 59974 26138
rect 60026 26086 60038 26138
rect 60090 26086 60102 26138
rect 60154 26086 89294 26138
rect 89346 26086 89358 26138
rect 89410 26086 89422 26138
rect 89474 26086 89486 26138
rect 89538 26086 89550 26138
rect 89602 26086 118864 26138
rect 1104 26064 118864 26086
rect 1394 26024 1400 26036
rect 1355 25996 1400 26024
rect 1394 25984 1400 25996
rect 1452 25984 1458 26036
rect 29086 25984 29092 26036
rect 29144 26024 29150 26036
rect 31662 26024 31668 26036
rect 29144 25996 31668 26024
rect 29144 25984 29150 25996
rect 31662 25984 31668 25996
rect 31720 25984 31726 26036
rect 31754 25984 31760 26036
rect 31812 26024 31818 26036
rect 34882 26024 34888 26036
rect 31812 25996 34888 26024
rect 31812 25984 31818 25996
rect 34882 25984 34888 25996
rect 34940 25984 34946 26036
rect 35253 26027 35311 26033
rect 35253 25993 35265 26027
rect 35299 26024 35311 26027
rect 36630 26024 36636 26036
rect 35299 25996 36636 26024
rect 35299 25993 35311 25996
rect 35253 25987 35311 25993
rect 36630 25984 36636 25996
rect 36688 25984 36694 26036
rect 50798 25984 50804 26036
rect 50856 26024 50862 26036
rect 55674 26024 55680 26036
rect 50856 25996 55680 26024
rect 50856 25984 50862 25996
rect 55674 25984 55680 25996
rect 55732 25984 55738 26036
rect 59909 26027 59967 26033
rect 59909 25993 59921 26027
rect 59955 26024 59967 26027
rect 60274 26024 60280 26036
rect 59955 25996 60280 26024
rect 59955 25993 59967 25996
rect 59909 25987 59967 25993
rect 60274 25984 60280 25996
rect 60332 25984 60338 26036
rect 61657 26027 61715 26033
rect 61657 25993 61669 26027
rect 61703 26024 61715 26027
rect 63310 26024 63316 26036
rect 61703 25996 63316 26024
rect 61703 25993 61715 25996
rect 61657 25987 61715 25993
rect 63310 25984 63316 25996
rect 63368 25984 63374 26036
rect 68554 25984 68560 26036
rect 68612 26024 68618 26036
rect 72050 26024 72056 26036
rect 68612 25996 72056 26024
rect 68612 25984 68618 25996
rect 72050 25984 72056 25996
rect 72108 25984 72114 26036
rect 76098 26024 76104 26036
rect 76059 25996 76104 26024
rect 76098 25984 76104 25996
rect 76156 25984 76162 26036
rect 77478 25984 77484 26036
rect 77536 26024 77542 26036
rect 85022 26024 85028 26036
rect 77536 25996 85028 26024
rect 77536 25984 77542 25996
rect 85022 25984 85028 25996
rect 85080 25984 85086 26036
rect 117225 26027 117283 26033
rect 117225 26024 117237 26027
rect 99346 25996 117237 26024
rect 54478 25956 54484 25968
rect 6886 25928 54484 25956
rect 1581 25891 1639 25897
rect 1581 25857 1593 25891
rect 1627 25888 1639 25891
rect 6886 25888 6914 25928
rect 54478 25916 54484 25928
rect 54536 25916 54542 25968
rect 58158 25956 58164 25968
rect 57900 25928 58164 25956
rect 1627 25860 6914 25888
rect 1627 25857 1639 25860
rect 1581 25851 1639 25857
rect 35250 25848 35256 25900
rect 35308 25888 35314 25900
rect 35437 25891 35495 25897
rect 35437 25888 35449 25891
rect 35308 25860 35449 25888
rect 35308 25848 35314 25860
rect 35437 25857 35449 25860
rect 35483 25857 35495 25891
rect 35437 25851 35495 25857
rect 40954 25848 40960 25900
rect 41012 25888 41018 25900
rect 46750 25888 46756 25900
rect 41012 25860 46756 25888
rect 41012 25848 41018 25860
rect 46750 25848 46756 25860
rect 46808 25848 46814 25900
rect 49970 25848 49976 25900
rect 50028 25888 50034 25900
rect 54110 25888 54116 25900
rect 50028 25860 54116 25888
rect 50028 25848 50034 25860
rect 54110 25848 54116 25860
rect 54168 25848 54174 25900
rect 57900 25897 57928 25928
rect 58158 25916 58164 25928
rect 58216 25956 58222 25968
rect 68278 25956 68284 25968
rect 58216 25928 68284 25956
rect 58216 25916 58222 25928
rect 68278 25916 68284 25928
rect 68336 25916 68342 25968
rect 71314 25916 71320 25968
rect 71372 25956 71378 25968
rect 81158 25956 81164 25968
rect 71372 25928 81164 25956
rect 71372 25916 71378 25928
rect 81158 25916 81164 25928
rect 81216 25916 81222 25968
rect 57885 25891 57943 25897
rect 57885 25857 57897 25891
rect 57931 25857 57943 25891
rect 57885 25851 57943 25857
rect 58066 25848 58072 25900
rect 58124 25888 58130 25900
rect 58526 25888 58532 25900
rect 58124 25860 58532 25888
rect 58124 25848 58130 25860
rect 58526 25848 58532 25860
rect 58584 25848 58590 25900
rect 60277 25891 60335 25897
rect 60277 25857 60289 25891
rect 60323 25857 60335 25891
rect 61838 25888 61844 25900
rect 61799 25860 61844 25888
rect 60277 25851 60335 25857
rect 56778 25780 56784 25832
rect 56836 25820 56842 25832
rect 60292 25820 60320 25851
rect 61838 25848 61844 25860
rect 61896 25848 61902 25900
rect 68002 25848 68008 25900
rect 68060 25888 68066 25900
rect 72786 25888 72792 25900
rect 68060 25860 72792 25888
rect 68060 25848 68066 25860
rect 72786 25848 72792 25860
rect 72844 25848 72850 25900
rect 76282 25888 76288 25900
rect 76243 25860 76288 25888
rect 76282 25848 76288 25860
rect 76340 25848 76346 25900
rect 77570 25848 77576 25900
rect 77628 25888 77634 25900
rect 82262 25888 82268 25900
rect 77628 25860 82268 25888
rect 77628 25848 77634 25860
rect 82262 25848 82268 25860
rect 82320 25848 82326 25900
rect 56836 25792 60320 25820
rect 56836 25780 56842 25792
rect 60366 25780 60372 25832
rect 60424 25820 60430 25832
rect 60553 25823 60611 25829
rect 60424 25792 60469 25820
rect 60424 25780 60430 25792
rect 60553 25789 60565 25823
rect 60599 25820 60611 25823
rect 64138 25820 64144 25832
rect 60599 25792 64144 25820
rect 60599 25789 60611 25792
rect 60553 25783 60611 25789
rect 64138 25780 64144 25792
rect 64196 25780 64202 25832
rect 76834 25820 76840 25832
rect 70366 25792 76840 25820
rect 60918 25752 60924 25764
rect 58544 25724 60924 25752
rect 58544 25696 58572 25724
rect 60918 25712 60924 25724
rect 60976 25712 60982 25764
rect 61010 25712 61016 25764
rect 61068 25752 61074 25764
rect 70366 25752 70394 25792
rect 76834 25780 76840 25792
rect 76892 25780 76898 25832
rect 61068 25724 70394 25752
rect 61068 25712 61074 25724
rect 94682 25712 94688 25764
rect 94740 25752 94746 25764
rect 99346 25752 99374 25996
rect 117225 25993 117237 25996
rect 117271 25993 117283 26027
rect 117225 25987 117283 25993
rect 117961 25959 118019 25965
rect 117961 25925 117973 25959
rect 118007 25956 118019 25959
rect 119798 25956 119804 25968
rect 118007 25928 119804 25956
rect 118007 25925 118019 25928
rect 117961 25919 118019 25925
rect 119798 25916 119804 25928
rect 119856 25916 119862 25968
rect 117409 25891 117467 25897
rect 117409 25857 117421 25891
rect 117455 25888 117467 25891
rect 117866 25888 117872 25900
rect 117455 25860 117872 25888
rect 117455 25857 117467 25860
rect 117409 25851 117467 25857
rect 117866 25848 117872 25860
rect 117924 25848 117930 25900
rect 118145 25755 118203 25761
rect 118145 25752 118157 25755
rect 94740 25724 99374 25752
rect 113744 25724 118157 25752
rect 94740 25712 94746 25724
rect 57882 25644 57888 25696
rect 57940 25684 57946 25696
rect 58253 25687 58311 25693
rect 58253 25684 58265 25687
rect 57940 25656 58265 25684
rect 57940 25644 57946 25656
rect 58253 25653 58265 25656
rect 58299 25653 58311 25687
rect 58526 25684 58532 25696
rect 58487 25656 58532 25684
rect 58253 25647 58311 25653
rect 58526 25644 58532 25656
rect 58584 25644 58590 25696
rect 59446 25644 59452 25696
rect 59504 25684 59510 25696
rect 59541 25687 59599 25693
rect 59541 25684 59553 25687
rect 59504 25656 59553 25684
rect 59504 25644 59510 25656
rect 59541 25653 59553 25656
rect 59587 25684 59599 25687
rect 60366 25684 60372 25696
rect 59587 25656 60372 25684
rect 59587 25653 59599 25656
rect 59541 25647 59599 25653
rect 60366 25644 60372 25656
rect 60424 25644 60430 25696
rect 78858 25644 78864 25696
rect 78916 25684 78922 25696
rect 113744 25684 113772 25724
rect 118145 25721 118157 25724
rect 118191 25721 118203 25755
rect 118145 25715 118203 25721
rect 78916 25656 113772 25684
rect 78916 25644 78922 25656
rect 1104 25594 118864 25616
rect 1104 25542 15674 25594
rect 15726 25542 15738 25594
rect 15790 25542 15802 25594
rect 15854 25542 15866 25594
rect 15918 25542 15930 25594
rect 15982 25542 45122 25594
rect 45174 25542 45186 25594
rect 45238 25542 45250 25594
rect 45302 25542 45314 25594
rect 45366 25542 45378 25594
rect 45430 25542 74570 25594
rect 74622 25542 74634 25594
rect 74686 25542 74698 25594
rect 74750 25542 74762 25594
rect 74814 25542 74826 25594
rect 74878 25542 104018 25594
rect 104070 25542 104082 25594
rect 104134 25542 104146 25594
rect 104198 25542 104210 25594
rect 104262 25542 104274 25594
rect 104326 25542 118864 25594
rect 1104 25520 118864 25542
rect 4430 25440 4436 25492
rect 4488 25480 4494 25492
rect 59446 25480 59452 25492
rect 4488 25452 59452 25480
rect 4488 25440 4494 25452
rect 59446 25440 59452 25452
rect 59504 25440 59510 25492
rect 32677 25415 32735 25421
rect 32677 25381 32689 25415
rect 32723 25412 32735 25415
rect 45097 25415 45155 25421
rect 32723 25384 41414 25412
rect 32723 25381 32735 25384
rect 32677 25375 32735 25381
rect 41386 25344 41414 25384
rect 45097 25381 45109 25415
rect 45143 25412 45155 25415
rect 45143 25384 51074 25412
rect 45143 25381 45155 25384
rect 45097 25375 45155 25381
rect 47210 25344 47216 25356
rect 41386 25316 47216 25344
rect 47210 25304 47216 25316
rect 47268 25304 47274 25356
rect 51046 25344 51074 25384
rect 54478 25372 54484 25424
rect 54536 25412 54542 25424
rect 58069 25415 58127 25421
rect 58069 25412 58081 25415
rect 54536 25384 58081 25412
rect 54536 25372 54542 25384
rect 58069 25381 58081 25384
rect 58115 25381 58127 25415
rect 58069 25375 58127 25381
rect 56870 25344 56876 25356
rect 51046 25316 56876 25344
rect 56870 25304 56876 25316
rect 56928 25304 56934 25356
rect 32858 25276 32864 25288
rect 32819 25248 32864 25276
rect 32858 25236 32864 25248
rect 32916 25236 32922 25288
rect 42702 25236 42708 25288
rect 42760 25276 42766 25288
rect 45281 25279 45339 25285
rect 45281 25276 45293 25279
rect 42760 25248 45293 25276
rect 42760 25236 42766 25248
rect 45281 25245 45293 25248
rect 45327 25245 45339 25279
rect 57882 25276 57888 25288
rect 57843 25248 57888 25276
rect 45281 25239 45339 25245
rect 57882 25236 57888 25248
rect 57940 25236 57946 25288
rect 64046 25276 64052 25288
rect 64007 25248 64052 25276
rect 64046 25236 64052 25248
rect 64104 25236 64110 25288
rect 107654 25236 107660 25288
rect 107712 25276 107718 25288
rect 118145 25279 118203 25285
rect 118145 25276 118157 25279
rect 107712 25248 118157 25276
rect 107712 25236 107718 25248
rect 118145 25245 118157 25248
rect 118191 25245 118203 25279
rect 118145 25239 118203 25245
rect 34514 25168 34520 25220
rect 34572 25208 34578 25220
rect 36633 25211 36691 25217
rect 36633 25208 36645 25211
rect 34572 25180 36645 25208
rect 34572 25168 34578 25180
rect 36633 25177 36645 25180
rect 36679 25177 36691 25211
rect 36633 25171 36691 25177
rect 36817 25211 36875 25217
rect 36817 25177 36829 25211
rect 36863 25208 36875 25211
rect 64230 25208 64236 25220
rect 36863 25180 60734 25208
rect 64191 25180 64236 25208
rect 36863 25177 36875 25180
rect 36817 25171 36875 25177
rect 60706 25140 60734 25180
rect 64230 25168 64236 25180
rect 64288 25168 64294 25220
rect 86402 25140 86408 25152
rect 60706 25112 86408 25140
rect 86402 25100 86408 25112
rect 86460 25100 86466 25152
rect 117958 25140 117964 25152
rect 117919 25112 117964 25140
rect 117958 25100 117964 25112
rect 118016 25100 118022 25152
rect 1104 25050 118864 25072
rect 1104 24998 30398 25050
rect 30450 24998 30462 25050
rect 30514 24998 30526 25050
rect 30578 24998 30590 25050
rect 30642 24998 30654 25050
rect 30706 24998 59846 25050
rect 59898 24998 59910 25050
rect 59962 24998 59974 25050
rect 60026 24998 60038 25050
rect 60090 24998 60102 25050
rect 60154 24998 89294 25050
rect 89346 24998 89358 25050
rect 89410 24998 89422 25050
rect 89474 24998 89486 25050
rect 89538 24998 89550 25050
rect 89602 24998 118864 25050
rect 1104 24976 118864 24998
rect 29546 24896 29552 24948
rect 29604 24936 29610 24948
rect 31021 24939 31079 24945
rect 31021 24936 31033 24939
rect 29604 24908 31033 24936
rect 29604 24896 29610 24908
rect 31021 24905 31033 24908
rect 31067 24905 31079 24939
rect 31021 24899 31079 24905
rect 32125 24939 32183 24945
rect 32125 24905 32137 24939
rect 32171 24936 32183 24939
rect 32858 24936 32864 24948
rect 32171 24908 32864 24936
rect 32171 24905 32183 24908
rect 32125 24899 32183 24905
rect 32858 24896 32864 24908
rect 32916 24896 32922 24948
rect 30944 24840 31156 24868
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24800 1731 24803
rect 30944 24800 30972 24840
rect 1719 24772 30972 24800
rect 31128 24800 31156 24840
rect 31128 24772 31432 24800
rect 1719 24769 1731 24772
rect 1673 24763 1731 24769
rect 1394 24732 1400 24744
rect 1355 24704 1400 24732
rect 1394 24692 1400 24704
rect 1452 24692 1458 24744
rect 31110 24732 31116 24744
rect 31071 24704 31116 24732
rect 31110 24692 31116 24704
rect 31168 24692 31174 24744
rect 31294 24732 31300 24744
rect 31255 24704 31300 24732
rect 31294 24692 31300 24704
rect 31352 24692 31358 24744
rect 31404 24732 31432 24772
rect 31754 24760 31760 24812
rect 31812 24800 31818 24812
rect 32493 24803 32551 24809
rect 32493 24800 32505 24803
rect 31812 24772 32505 24800
rect 31812 24760 31818 24772
rect 32493 24769 32505 24772
rect 32539 24769 32551 24803
rect 118145 24803 118203 24809
rect 118145 24800 118157 24803
rect 32493 24763 32551 24769
rect 117608 24772 118157 24800
rect 32585 24735 32643 24741
rect 32585 24732 32597 24735
rect 31404 24704 32597 24732
rect 32585 24701 32597 24704
rect 32631 24701 32643 24735
rect 32585 24695 32643 24701
rect 32769 24735 32827 24741
rect 32769 24701 32781 24735
rect 32815 24732 32827 24735
rect 32858 24732 32864 24744
rect 32815 24704 32864 24732
rect 32815 24701 32827 24704
rect 32769 24695 32827 24701
rect 32858 24692 32864 24704
rect 32916 24732 32922 24744
rect 33229 24735 33287 24741
rect 33229 24732 33241 24735
rect 32916 24704 33241 24732
rect 32916 24692 32922 24704
rect 33229 24701 33241 24704
rect 33275 24732 33287 24735
rect 33275 24704 51074 24732
rect 33275 24701 33287 24704
rect 33229 24695 33287 24701
rect 30653 24667 30711 24673
rect 30653 24633 30665 24667
rect 30699 24664 30711 24667
rect 42702 24664 42708 24676
rect 30699 24636 42708 24664
rect 30699 24633 30711 24636
rect 30653 24627 30711 24633
rect 42702 24624 42708 24636
rect 42760 24624 42766 24676
rect 31754 24556 31760 24608
rect 31812 24596 31818 24608
rect 51046 24596 51074 24704
rect 59630 24596 59636 24608
rect 31812 24568 31857 24596
rect 51046 24568 59636 24596
rect 31812 24556 31818 24568
rect 59630 24556 59636 24568
rect 59688 24556 59694 24608
rect 64230 24556 64236 24608
rect 64288 24596 64294 24608
rect 117608 24605 117636 24772
rect 118145 24769 118157 24772
rect 118191 24769 118203 24803
rect 118145 24763 118203 24769
rect 117593 24599 117651 24605
rect 117593 24596 117605 24599
rect 64288 24568 117605 24596
rect 64288 24556 64294 24568
rect 117593 24565 117605 24568
rect 117639 24565 117651 24599
rect 117958 24596 117964 24608
rect 117919 24568 117964 24596
rect 117593 24559 117651 24565
rect 117958 24556 117964 24568
rect 118016 24556 118022 24608
rect 1104 24506 118864 24528
rect 1104 24454 15674 24506
rect 15726 24454 15738 24506
rect 15790 24454 15802 24506
rect 15854 24454 15866 24506
rect 15918 24454 15930 24506
rect 15982 24454 45122 24506
rect 45174 24454 45186 24506
rect 45238 24454 45250 24506
rect 45302 24454 45314 24506
rect 45366 24454 45378 24506
rect 45430 24454 74570 24506
rect 74622 24454 74634 24506
rect 74686 24454 74698 24506
rect 74750 24454 74762 24506
rect 74814 24454 74826 24506
rect 74878 24454 104018 24506
rect 104070 24454 104082 24506
rect 104134 24454 104146 24506
rect 104198 24454 104210 24506
rect 104262 24454 104274 24506
rect 104326 24454 118864 24506
rect 1104 24432 118864 24454
rect 30653 24395 30711 24401
rect 30653 24361 30665 24395
rect 30699 24392 30711 24395
rect 34514 24392 34520 24404
rect 30699 24364 34520 24392
rect 30699 24361 30711 24364
rect 30653 24355 30711 24361
rect 34514 24352 34520 24364
rect 34572 24352 34578 24404
rect 31294 24256 31300 24268
rect 31255 24228 31300 24256
rect 31294 24216 31300 24228
rect 31352 24216 31358 24268
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24148 1458 24200
rect 1670 24188 1676 24200
rect 1631 24160 1676 24188
rect 1670 24148 1676 24160
rect 1728 24148 1734 24200
rect 2682 24148 2688 24200
rect 2740 24148 2746 24200
rect 2869 24191 2927 24197
rect 2869 24157 2881 24191
rect 2915 24188 2927 24191
rect 2958 24188 2964 24200
rect 2915 24160 2964 24188
rect 2915 24157 2927 24160
rect 2869 24151 2927 24157
rect 2958 24148 2964 24160
rect 3016 24148 3022 24200
rect 51074 24148 51080 24200
rect 51132 24188 51138 24200
rect 51442 24188 51448 24200
rect 51132 24160 51448 24188
rect 51132 24148 51138 24160
rect 51442 24148 51448 24160
rect 51500 24148 51506 24200
rect 2700 24120 2728 24148
rect 30377 24123 30435 24129
rect 30377 24120 30389 24123
rect 2700 24092 30389 24120
rect 30377 24089 30389 24092
rect 30423 24120 30435 24123
rect 31021 24123 31079 24129
rect 31021 24120 31033 24123
rect 30423 24092 31033 24120
rect 30423 24089 30435 24092
rect 30377 24083 30435 24089
rect 31021 24089 31033 24092
rect 31067 24089 31079 24123
rect 31021 24083 31079 24089
rect 35434 24080 35440 24132
rect 35492 24120 35498 24132
rect 102226 24120 102232 24132
rect 35492 24092 102232 24120
rect 35492 24080 35498 24092
rect 102226 24080 102232 24092
rect 102284 24080 102290 24132
rect 1486 24012 1492 24064
rect 1544 24052 1550 24064
rect 2685 24055 2743 24061
rect 2685 24052 2697 24055
rect 1544 24024 2697 24052
rect 1544 24012 1550 24024
rect 2685 24021 2697 24024
rect 2731 24021 2743 24055
rect 2685 24015 2743 24021
rect 28810 24012 28816 24064
rect 28868 24052 28874 24064
rect 31113 24055 31171 24061
rect 31113 24052 31125 24055
rect 28868 24024 31125 24052
rect 28868 24012 28874 24024
rect 31113 24021 31125 24024
rect 31159 24021 31171 24055
rect 31113 24015 31171 24021
rect 1104 23962 118864 23984
rect 1104 23910 30398 23962
rect 30450 23910 30462 23962
rect 30514 23910 30526 23962
rect 30578 23910 30590 23962
rect 30642 23910 30654 23962
rect 30706 23910 59846 23962
rect 59898 23910 59910 23962
rect 59962 23910 59974 23962
rect 60026 23910 60038 23962
rect 60090 23910 60102 23962
rect 60154 23910 89294 23962
rect 89346 23910 89358 23962
rect 89410 23910 89422 23962
rect 89474 23910 89486 23962
rect 89538 23910 89550 23962
rect 89602 23910 118864 23962
rect 1104 23888 118864 23910
rect 1581 23715 1639 23721
rect 1581 23681 1593 23715
rect 1627 23712 1639 23715
rect 1762 23712 1768 23724
rect 1627 23684 1768 23712
rect 1627 23681 1639 23684
rect 1581 23675 1639 23681
rect 1762 23672 1768 23684
rect 1820 23672 1826 23724
rect 91002 23672 91008 23724
rect 91060 23712 91066 23724
rect 117593 23715 117651 23721
rect 117593 23712 117605 23715
rect 91060 23684 117605 23712
rect 91060 23672 91066 23684
rect 117593 23681 117605 23684
rect 117639 23681 117651 23715
rect 117593 23675 117651 23681
rect 117222 23604 117228 23656
rect 117280 23644 117286 23656
rect 117317 23647 117375 23653
rect 117317 23644 117329 23647
rect 117280 23616 117329 23644
rect 117280 23604 117286 23616
rect 117317 23613 117329 23616
rect 117363 23613 117375 23647
rect 117317 23607 117375 23613
rect 1394 23508 1400 23520
rect 1355 23480 1400 23508
rect 1394 23468 1400 23480
rect 1452 23468 1458 23520
rect 1104 23418 118864 23440
rect 1104 23366 15674 23418
rect 15726 23366 15738 23418
rect 15790 23366 15802 23418
rect 15854 23366 15866 23418
rect 15918 23366 15930 23418
rect 15982 23366 45122 23418
rect 45174 23366 45186 23418
rect 45238 23366 45250 23418
rect 45302 23366 45314 23418
rect 45366 23366 45378 23418
rect 45430 23366 74570 23418
rect 74622 23366 74634 23418
rect 74686 23366 74698 23418
rect 74750 23366 74762 23418
rect 74814 23366 74826 23418
rect 74878 23366 104018 23418
rect 104070 23366 104082 23418
rect 104134 23366 104146 23418
rect 104198 23366 104210 23418
rect 104262 23366 104274 23418
rect 104326 23366 118864 23418
rect 1104 23344 118864 23366
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 11698 22964 11704 22976
rect 1728 22936 11704 22964
rect 1728 22924 1734 22936
rect 11698 22924 11704 22936
rect 11756 22924 11762 22976
rect 14642 22924 14648 22976
rect 14700 22964 14706 22976
rect 71222 22964 71228 22976
rect 14700 22936 71228 22964
rect 14700 22924 14706 22936
rect 71222 22924 71228 22936
rect 71280 22924 71286 22976
rect 1104 22874 118864 22896
rect 1104 22822 30398 22874
rect 30450 22822 30462 22874
rect 30514 22822 30526 22874
rect 30578 22822 30590 22874
rect 30642 22822 30654 22874
rect 30706 22822 59846 22874
rect 59898 22822 59910 22874
rect 59962 22822 59974 22874
rect 60026 22822 60038 22874
rect 60090 22822 60102 22874
rect 60154 22822 89294 22874
rect 89346 22822 89358 22874
rect 89410 22822 89422 22874
rect 89474 22822 89486 22874
rect 89538 22822 89550 22874
rect 89602 22822 118864 22874
rect 1104 22800 118864 22822
rect 9214 22720 9220 22772
rect 9272 22760 9278 22772
rect 98178 22760 98184 22772
rect 9272 22732 98184 22760
rect 9272 22720 9278 22732
rect 98178 22720 98184 22732
rect 98236 22720 98242 22772
rect 88794 22652 88800 22704
rect 88852 22692 88858 22704
rect 94869 22695 94927 22701
rect 94869 22692 94881 22695
rect 88852 22664 94881 22692
rect 88852 22652 88858 22664
rect 94869 22661 94881 22664
rect 94915 22661 94927 22695
rect 94869 22655 94927 22661
rect 94774 22624 94780 22636
rect 94735 22596 94780 22624
rect 94774 22584 94780 22596
rect 94832 22584 94838 22636
rect 95789 22627 95847 22633
rect 95789 22593 95801 22627
rect 95835 22593 95847 22627
rect 118145 22627 118203 22633
rect 118145 22624 118157 22627
rect 95789 22587 95847 22593
rect 99346 22596 118157 22624
rect 94958 22556 94964 22568
rect 94919 22528 94964 22556
rect 94958 22516 94964 22528
rect 95016 22556 95022 22568
rect 95421 22559 95479 22565
rect 95421 22556 95433 22559
rect 95016 22528 95433 22556
rect 95016 22516 95022 22528
rect 95421 22525 95433 22528
rect 95467 22525 95479 22559
rect 95421 22519 95479 22525
rect 94409 22491 94467 22497
rect 94409 22457 94421 22491
rect 94455 22488 94467 22491
rect 95804 22488 95832 22587
rect 94455 22460 95832 22488
rect 94455 22457 94467 22460
rect 94409 22451 94467 22457
rect 95605 22423 95663 22429
rect 95605 22389 95617 22423
rect 95651 22420 95663 22423
rect 99346 22420 99374 22596
rect 118145 22593 118157 22596
rect 118191 22593 118203 22627
rect 118145 22587 118203 22593
rect 117958 22488 117964 22500
rect 117919 22460 117964 22488
rect 117958 22448 117964 22460
rect 118016 22448 118022 22500
rect 95651 22392 99374 22420
rect 95651 22389 95663 22392
rect 95605 22383 95663 22389
rect 1104 22330 118864 22352
rect 1104 22278 15674 22330
rect 15726 22278 15738 22330
rect 15790 22278 15802 22330
rect 15854 22278 15866 22330
rect 15918 22278 15930 22330
rect 15982 22278 45122 22330
rect 45174 22278 45186 22330
rect 45238 22278 45250 22330
rect 45302 22278 45314 22330
rect 45366 22278 45378 22330
rect 45430 22278 74570 22330
rect 74622 22278 74634 22330
rect 74686 22278 74698 22330
rect 74750 22278 74762 22330
rect 74814 22278 74826 22330
rect 74878 22278 104018 22330
rect 104070 22278 104082 22330
rect 104134 22278 104146 22330
rect 104198 22278 104210 22330
rect 104262 22278 104274 22330
rect 104326 22278 118864 22330
rect 1104 22256 118864 22278
rect 50706 22080 50712 22092
rect 50667 22052 50712 22080
rect 50706 22040 50712 22052
rect 50764 22040 50770 22092
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 22012 1639 22015
rect 49513 22015 49571 22021
rect 49513 22012 49525 22015
rect 1627 21984 49525 22012
rect 1627 21981 1639 21984
rect 1581 21975 1639 21981
rect 49513 21981 49525 21984
rect 49559 21981 49571 22015
rect 49513 21975 49571 21981
rect 50525 22015 50583 22021
rect 50525 21981 50537 22015
rect 50571 22012 50583 22015
rect 51074 22012 51080 22024
rect 50571 21984 51080 22012
rect 50571 21981 50583 21984
rect 50525 21975 50583 21981
rect 51074 21972 51080 21984
rect 51132 21972 51138 22024
rect 49329 21947 49387 21953
rect 49329 21913 49341 21947
rect 49375 21944 49387 21947
rect 49375 21916 50200 21944
rect 49375 21913 49387 21916
rect 49329 21907 49387 21913
rect 1394 21876 1400 21888
rect 1355 21848 1400 21876
rect 1394 21836 1400 21848
rect 1452 21836 1458 21888
rect 50172 21885 50200 21916
rect 68186 21904 68192 21956
rect 68244 21944 68250 21956
rect 68557 21947 68615 21953
rect 68557 21944 68569 21947
rect 68244 21916 68569 21944
rect 68244 21904 68250 21916
rect 68557 21913 68569 21916
rect 68603 21913 68615 21947
rect 68557 21907 68615 21913
rect 50157 21879 50215 21885
rect 50157 21845 50169 21879
rect 50203 21845 50215 21879
rect 50157 21839 50215 21845
rect 50614 21836 50620 21888
rect 50672 21876 50678 21888
rect 68649 21879 68707 21885
rect 50672 21848 50717 21876
rect 50672 21836 50678 21848
rect 68649 21845 68661 21879
rect 68695 21876 68707 21879
rect 106366 21876 106372 21888
rect 68695 21848 106372 21876
rect 68695 21845 68707 21848
rect 68649 21839 68707 21845
rect 106366 21836 106372 21848
rect 106424 21836 106430 21888
rect 1104 21786 118864 21808
rect 1104 21734 30398 21786
rect 30450 21734 30462 21786
rect 30514 21734 30526 21786
rect 30578 21734 30590 21786
rect 30642 21734 30654 21786
rect 30706 21734 59846 21786
rect 59898 21734 59910 21786
rect 59962 21734 59974 21786
rect 60026 21734 60038 21786
rect 60090 21734 60102 21786
rect 60154 21734 89294 21786
rect 89346 21734 89358 21786
rect 89410 21734 89422 21786
rect 89474 21734 89486 21786
rect 89538 21734 89550 21786
rect 89602 21734 118864 21786
rect 1104 21712 118864 21734
rect 47765 21675 47823 21681
rect 47765 21641 47777 21675
rect 47811 21672 47823 21675
rect 49694 21672 49700 21684
rect 47811 21644 49700 21672
rect 47811 21641 47823 21644
rect 47765 21635 47823 21641
rect 49694 21632 49700 21644
rect 49752 21672 49758 21684
rect 50706 21672 50712 21684
rect 49752 21644 50712 21672
rect 49752 21632 49758 21644
rect 50706 21632 50712 21644
rect 50764 21632 50770 21684
rect 68186 21672 68192 21684
rect 68147 21644 68192 21672
rect 68186 21632 68192 21644
rect 68244 21632 68250 21684
rect 1394 21536 1400 21548
rect 1355 21508 1400 21536
rect 1394 21496 1400 21508
rect 1452 21496 1458 21548
rect 47581 21539 47639 21545
rect 47581 21505 47593 21539
rect 47627 21536 47639 21539
rect 54478 21536 54484 21548
rect 47627 21508 54484 21536
rect 47627 21505 47639 21508
rect 47581 21499 47639 21505
rect 54478 21496 54484 21508
rect 54536 21496 54542 21548
rect 68094 21496 68100 21548
rect 68152 21536 68158 21548
rect 68557 21539 68615 21545
rect 68557 21536 68569 21539
rect 68152 21508 68569 21536
rect 68152 21496 68158 21508
rect 68557 21505 68569 21508
rect 68603 21505 68615 21539
rect 68557 21499 68615 21505
rect 68646 21468 68652 21480
rect 68607 21440 68652 21468
rect 68646 21428 68652 21440
rect 68704 21428 68710 21480
rect 68738 21428 68744 21480
rect 68796 21468 68802 21480
rect 79226 21468 79232 21480
rect 68796 21440 79232 21468
rect 68796 21428 68802 21440
rect 79226 21428 79232 21440
rect 79284 21428 79290 21480
rect 117314 21468 117320 21480
rect 117275 21440 117320 21468
rect 117314 21428 117320 21440
rect 117372 21428 117378 21480
rect 117590 21468 117596 21480
rect 117551 21440 117596 21468
rect 117590 21428 117596 21440
rect 117648 21428 117654 21480
rect 28902 21360 28908 21412
rect 28960 21400 28966 21412
rect 82722 21400 82728 21412
rect 28960 21372 82728 21400
rect 28960 21360 28966 21372
rect 82722 21360 82728 21372
rect 82780 21360 82786 21412
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 1104 21242 118864 21264
rect 1104 21190 15674 21242
rect 15726 21190 15738 21242
rect 15790 21190 15802 21242
rect 15854 21190 15866 21242
rect 15918 21190 15930 21242
rect 15982 21190 45122 21242
rect 45174 21190 45186 21242
rect 45238 21190 45250 21242
rect 45302 21190 45314 21242
rect 45366 21190 45378 21242
rect 45430 21190 74570 21242
rect 74622 21190 74634 21242
rect 74686 21190 74698 21242
rect 74750 21190 74762 21242
rect 74814 21190 74826 21242
rect 74878 21190 104018 21242
rect 104070 21190 104082 21242
rect 104134 21190 104146 21242
rect 104198 21190 104210 21242
rect 104262 21190 104274 21242
rect 104326 21190 118864 21242
rect 1104 21168 118864 21190
rect 1578 21088 1584 21140
rect 1636 21128 1642 21140
rect 68646 21128 68652 21140
rect 1636 21100 68652 21128
rect 1636 21088 1642 21100
rect 68646 21088 68652 21100
rect 68704 21088 68710 21140
rect 54665 21063 54723 21069
rect 54665 21029 54677 21063
rect 54711 21060 54723 21063
rect 55122 21060 55128 21072
rect 54711 21032 55128 21060
rect 54711 21029 54723 21032
rect 54665 21023 54723 21029
rect 55122 21020 55128 21032
rect 55180 21020 55186 21072
rect 117590 21060 117596 21072
rect 84856 21032 117596 21060
rect 54570 20952 54576 21004
rect 54628 20992 54634 21004
rect 72878 20992 72884 21004
rect 54628 20964 56088 20992
rect 72839 20964 72884 20992
rect 54628 20952 54634 20964
rect 54478 20924 54484 20936
rect 54439 20896 54484 20924
rect 54478 20884 54484 20896
rect 54536 20924 54542 20936
rect 55490 20924 55496 20936
rect 54536 20896 55496 20924
rect 54536 20884 54542 20896
rect 55490 20884 55496 20896
rect 55548 20924 55554 20936
rect 55769 20927 55827 20933
rect 55769 20924 55781 20927
rect 55548 20896 55781 20924
rect 55548 20884 55554 20896
rect 55769 20893 55781 20896
rect 55815 20893 55827 20927
rect 55769 20887 55827 20893
rect 56060 20797 56088 20964
rect 72878 20952 72884 20964
rect 72936 20952 72942 21004
rect 72694 20924 72700 20936
rect 72655 20896 72700 20924
rect 72694 20884 72700 20896
rect 72752 20884 72758 20936
rect 84856 20933 84884 21032
rect 117590 21020 117596 21032
rect 117648 21020 117654 21072
rect 85022 20992 85028 21004
rect 84983 20964 85028 20992
rect 85022 20952 85028 20964
rect 85080 20952 85086 21004
rect 84841 20927 84899 20933
rect 84841 20893 84853 20927
rect 84887 20893 84899 20927
rect 84841 20887 84899 20893
rect 115934 20884 115940 20936
rect 115992 20924 115998 20936
rect 118145 20927 118203 20933
rect 118145 20924 118157 20927
rect 115992 20896 118157 20924
rect 115992 20884 115998 20896
rect 118145 20893 118157 20896
rect 118191 20893 118203 20927
rect 118145 20887 118203 20893
rect 84197 20859 84255 20865
rect 84197 20825 84209 20859
rect 84243 20856 84255 20859
rect 84933 20859 84991 20865
rect 84933 20856 84945 20859
rect 84243 20828 84945 20856
rect 84243 20825 84255 20828
rect 84197 20819 84255 20825
rect 84933 20825 84945 20828
rect 84979 20856 84991 20859
rect 118050 20856 118056 20868
rect 84979 20828 118056 20856
rect 84979 20825 84991 20828
rect 84933 20819 84991 20825
rect 118050 20816 118056 20828
rect 118108 20816 118114 20868
rect 56045 20791 56103 20797
rect 56045 20757 56057 20791
rect 56091 20788 56103 20791
rect 68738 20788 68744 20800
rect 56091 20760 68744 20788
rect 56091 20757 56103 20760
rect 56045 20751 56103 20757
rect 68738 20748 68744 20760
rect 68796 20748 68802 20800
rect 71866 20748 71872 20800
rect 71924 20788 71930 20800
rect 72329 20791 72387 20797
rect 72329 20788 72341 20791
rect 71924 20760 72341 20788
rect 71924 20748 71930 20760
rect 72329 20757 72341 20760
rect 72375 20757 72387 20791
rect 72329 20751 72387 20757
rect 72786 20748 72792 20800
rect 72844 20788 72850 20800
rect 84470 20788 84476 20800
rect 72844 20760 72889 20788
rect 84431 20760 84476 20788
rect 72844 20748 72850 20760
rect 84470 20748 84476 20760
rect 84528 20748 84534 20800
rect 117958 20788 117964 20800
rect 117919 20760 117964 20788
rect 117958 20748 117964 20760
rect 118016 20748 118022 20800
rect 1104 20698 118864 20720
rect 1104 20646 30398 20698
rect 30450 20646 30462 20698
rect 30514 20646 30526 20698
rect 30578 20646 30590 20698
rect 30642 20646 30654 20698
rect 30706 20646 59846 20698
rect 59898 20646 59910 20698
rect 59962 20646 59974 20698
rect 60026 20646 60038 20698
rect 60090 20646 60102 20698
rect 60154 20646 89294 20698
rect 89346 20646 89358 20698
rect 89410 20646 89422 20698
rect 89474 20646 89486 20698
rect 89538 20646 89550 20698
rect 89602 20646 118864 20698
rect 1104 20624 118864 20646
rect 79137 20587 79195 20593
rect 79137 20553 79149 20587
rect 79183 20584 79195 20587
rect 86862 20584 86868 20596
rect 79183 20556 86868 20584
rect 79183 20553 79195 20556
rect 79137 20547 79195 20553
rect 86862 20544 86868 20556
rect 86920 20544 86926 20596
rect 114557 20587 114615 20593
rect 114557 20553 114569 20587
rect 114603 20584 114615 20587
rect 115934 20584 115940 20596
rect 114603 20556 115940 20584
rect 114603 20553 114615 20556
rect 114557 20547 114615 20553
rect 115934 20544 115940 20556
rect 115992 20544 115998 20596
rect 71866 20448 71872 20460
rect 71827 20420 71872 20448
rect 71866 20408 71872 20420
rect 71924 20408 71930 20460
rect 79042 20448 79048 20460
rect 79003 20420 79048 20448
rect 79042 20408 79048 20420
rect 79100 20448 79106 20460
rect 79689 20451 79747 20457
rect 79689 20448 79701 20451
rect 79100 20420 79701 20448
rect 79100 20408 79106 20420
rect 79689 20417 79701 20420
rect 79735 20417 79747 20451
rect 79689 20411 79747 20417
rect 83645 20451 83703 20457
rect 83645 20417 83657 20451
rect 83691 20448 83703 20451
rect 84470 20448 84476 20460
rect 83691 20420 84476 20448
rect 83691 20417 83703 20420
rect 83645 20411 83703 20417
rect 84470 20408 84476 20420
rect 84528 20408 84534 20460
rect 114738 20448 114744 20460
rect 114699 20420 114744 20448
rect 114738 20408 114744 20420
rect 114796 20408 114802 20460
rect 79226 20380 79232 20392
rect 79187 20352 79232 20380
rect 79226 20340 79232 20352
rect 79284 20340 79290 20392
rect 83921 20383 83979 20389
rect 83921 20349 83933 20383
rect 83967 20349 83979 20383
rect 83921 20343 83979 20349
rect 78030 20272 78036 20324
rect 78088 20312 78094 20324
rect 83936 20312 83964 20343
rect 78088 20284 83964 20312
rect 78088 20272 78094 20284
rect 72050 20244 72056 20256
rect 72011 20216 72056 20244
rect 72050 20204 72056 20216
rect 72108 20204 72114 20256
rect 78674 20244 78680 20256
rect 78635 20216 78680 20244
rect 78674 20204 78680 20216
rect 78732 20204 78738 20256
rect 1104 20154 118864 20176
rect 1104 20102 15674 20154
rect 15726 20102 15738 20154
rect 15790 20102 15802 20154
rect 15854 20102 15866 20154
rect 15918 20102 15930 20154
rect 15982 20102 45122 20154
rect 45174 20102 45186 20154
rect 45238 20102 45250 20154
rect 45302 20102 45314 20154
rect 45366 20102 45378 20154
rect 45430 20102 74570 20154
rect 74622 20102 74634 20154
rect 74686 20102 74698 20154
rect 74750 20102 74762 20154
rect 74814 20102 74826 20154
rect 74878 20102 104018 20154
rect 104070 20102 104082 20154
rect 104134 20102 104146 20154
rect 104198 20102 104210 20154
rect 104262 20102 104274 20154
rect 104326 20102 118864 20154
rect 1104 20080 118864 20102
rect 47026 20000 47032 20052
rect 47084 20040 47090 20052
rect 79042 20040 79048 20052
rect 47084 20012 79048 20040
rect 47084 20000 47090 20012
rect 79042 20000 79048 20012
rect 79100 20000 79106 20052
rect 1581 19839 1639 19845
rect 1581 19805 1593 19839
rect 1627 19836 1639 19839
rect 72050 19836 72056 19848
rect 1627 19808 72056 19836
rect 1627 19805 1639 19808
rect 1581 19799 1639 19805
rect 72050 19796 72056 19808
rect 72108 19796 72114 19848
rect 78674 19796 78680 19848
rect 78732 19836 78738 19848
rect 80149 19839 80207 19845
rect 80149 19836 80161 19839
rect 78732 19808 80161 19836
rect 78732 19796 78738 19808
rect 80149 19805 80161 19808
rect 80195 19805 80207 19839
rect 118145 19839 118203 19845
rect 118145 19836 118157 19839
rect 80149 19799 80207 19805
rect 84166 19808 118157 19836
rect 78950 19728 78956 19780
rect 79008 19768 79014 19780
rect 79321 19771 79379 19777
rect 79321 19768 79333 19771
rect 79008 19740 79333 19768
rect 79008 19728 79014 19740
rect 79321 19737 79333 19740
rect 79367 19737 79379 19771
rect 79321 19731 79379 19737
rect 79505 19771 79563 19777
rect 79505 19737 79517 19771
rect 79551 19768 79563 19771
rect 84166 19768 84194 19808
rect 118145 19805 118157 19808
rect 118191 19805 118203 19839
rect 118145 19799 118203 19805
rect 79551 19740 84194 19768
rect 113637 19771 113695 19777
rect 79551 19737 79563 19740
rect 79505 19731 79563 19737
rect 113637 19737 113649 19771
rect 113683 19768 113695 19771
rect 114738 19768 114744 19780
rect 113683 19740 114744 19768
rect 113683 19737 113695 19740
rect 113637 19731 113695 19737
rect 114738 19728 114744 19740
rect 114796 19728 114802 19780
rect 1394 19700 1400 19712
rect 1355 19672 1400 19700
rect 1394 19660 1400 19672
rect 1452 19660 1458 19712
rect 79965 19703 80023 19709
rect 79965 19669 79977 19703
rect 80011 19700 80023 19703
rect 80698 19700 80704 19712
rect 80011 19672 80704 19700
rect 80011 19669 80023 19672
rect 79965 19663 80023 19669
rect 80698 19660 80704 19672
rect 80756 19660 80762 19712
rect 113726 19700 113732 19712
rect 113687 19672 113732 19700
rect 113726 19660 113732 19672
rect 113784 19660 113790 19712
rect 117958 19700 117964 19712
rect 117919 19672 117964 19700
rect 117958 19660 117964 19672
rect 118016 19660 118022 19712
rect 1104 19610 118864 19632
rect 1104 19558 30398 19610
rect 30450 19558 30462 19610
rect 30514 19558 30526 19610
rect 30578 19558 30590 19610
rect 30642 19558 30654 19610
rect 30706 19558 59846 19610
rect 59898 19558 59910 19610
rect 59962 19558 59974 19610
rect 60026 19558 60038 19610
rect 60090 19558 60102 19610
rect 60154 19558 89294 19610
rect 89346 19558 89358 19610
rect 89410 19558 89422 19610
rect 89474 19558 89486 19610
rect 89538 19558 89550 19610
rect 89602 19558 118864 19610
rect 1104 19536 118864 19558
rect 102686 19456 102692 19508
rect 102744 19496 102750 19508
rect 113726 19496 113732 19508
rect 102744 19468 113732 19496
rect 102744 19456 102750 19468
rect 113726 19456 113732 19468
rect 113784 19456 113790 19508
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 2133 19159 2191 19165
rect 2133 19125 2145 19159
rect 2179 19156 2191 19159
rect 66530 19156 66536 19168
rect 2179 19128 66536 19156
rect 2179 19125 2191 19128
rect 2133 19119 2191 19125
rect 66530 19116 66536 19128
rect 66588 19116 66594 19168
rect 1104 19066 118864 19088
rect 1104 19014 15674 19066
rect 15726 19014 15738 19066
rect 15790 19014 15802 19066
rect 15854 19014 15866 19066
rect 15918 19014 15930 19066
rect 15982 19014 45122 19066
rect 45174 19014 45186 19066
rect 45238 19014 45250 19066
rect 45302 19014 45314 19066
rect 45366 19014 45378 19066
rect 45430 19014 74570 19066
rect 74622 19014 74634 19066
rect 74686 19014 74698 19066
rect 74750 19014 74762 19066
rect 74814 19014 74826 19066
rect 74878 19014 104018 19066
rect 104070 19014 104082 19066
rect 104134 19014 104146 19066
rect 104198 19014 104210 19066
rect 104262 19014 104274 19066
rect 104326 19014 118864 19066
rect 1104 18992 118864 19014
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 33318 18748 33324 18760
rect 1627 18720 33324 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 33318 18708 33324 18720
rect 33376 18708 33382 18760
rect 117866 18748 117872 18760
rect 117827 18720 117872 18748
rect 117866 18708 117872 18720
rect 117924 18708 117930 18760
rect 2222 18640 2228 18692
rect 2280 18680 2286 18692
rect 68554 18680 68560 18692
rect 2280 18652 68560 18680
rect 2280 18640 2286 18652
rect 68554 18640 68560 18652
rect 68612 18640 68618 18692
rect 1394 18612 1400 18624
rect 1355 18584 1400 18612
rect 1394 18572 1400 18584
rect 1452 18572 1458 18624
rect 117958 18572 117964 18624
rect 118016 18612 118022 18624
rect 118053 18615 118111 18621
rect 118053 18612 118065 18615
rect 118016 18584 118065 18612
rect 118016 18572 118022 18584
rect 118053 18581 118065 18584
rect 118099 18581 118111 18615
rect 118053 18575 118111 18581
rect 1104 18522 118864 18544
rect 1104 18470 30398 18522
rect 30450 18470 30462 18522
rect 30514 18470 30526 18522
rect 30578 18470 30590 18522
rect 30642 18470 30654 18522
rect 30706 18470 59846 18522
rect 59898 18470 59910 18522
rect 59962 18470 59974 18522
rect 60026 18470 60038 18522
rect 60090 18470 60102 18522
rect 60154 18470 89294 18522
rect 89346 18470 89358 18522
rect 89410 18470 89422 18522
rect 89474 18470 89486 18522
rect 89538 18470 89550 18522
rect 89602 18470 118864 18522
rect 1104 18448 118864 18470
rect 33318 18272 33324 18284
rect 33279 18244 33324 18272
rect 33318 18232 33324 18244
rect 33376 18232 33382 18284
rect 117866 18272 117872 18284
rect 117827 18244 117872 18272
rect 117866 18232 117872 18244
rect 117924 18232 117930 18284
rect 33045 18207 33103 18213
rect 33045 18173 33057 18207
rect 33091 18204 33103 18207
rect 33226 18204 33232 18216
rect 33091 18176 33232 18204
rect 33091 18173 33103 18176
rect 33045 18167 33103 18173
rect 33226 18164 33232 18176
rect 33284 18164 33290 18216
rect 117682 18028 117688 18080
rect 117740 18068 117746 18080
rect 118053 18071 118111 18077
rect 118053 18068 118065 18071
rect 117740 18040 118065 18068
rect 117740 18028 117746 18040
rect 118053 18037 118065 18040
rect 118099 18037 118111 18071
rect 118053 18031 118111 18037
rect 1104 17978 118864 18000
rect 1104 17926 15674 17978
rect 15726 17926 15738 17978
rect 15790 17926 15802 17978
rect 15854 17926 15866 17978
rect 15918 17926 15930 17978
rect 15982 17926 45122 17978
rect 45174 17926 45186 17978
rect 45238 17926 45250 17978
rect 45302 17926 45314 17978
rect 45366 17926 45378 17978
rect 45430 17926 74570 17978
rect 74622 17926 74634 17978
rect 74686 17926 74698 17978
rect 74750 17926 74762 17978
rect 74814 17926 74826 17978
rect 74878 17926 104018 17978
rect 104070 17926 104082 17978
rect 104134 17926 104146 17978
rect 104198 17926 104210 17978
rect 104262 17926 104274 17978
rect 104326 17926 118864 17978
rect 1104 17904 118864 17926
rect 33226 17824 33232 17876
rect 33284 17864 33290 17876
rect 33321 17867 33379 17873
rect 33321 17864 33333 17867
rect 33284 17836 33333 17864
rect 33284 17824 33290 17836
rect 33321 17833 33333 17836
rect 33367 17833 33379 17867
rect 33321 17827 33379 17833
rect 81434 17756 81440 17808
rect 81492 17796 81498 17808
rect 82722 17796 82728 17808
rect 81492 17768 82728 17796
rect 81492 17756 81498 17768
rect 82722 17756 82728 17768
rect 82780 17756 82786 17808
rect 31294 17688 31300 17740
rect 31352 17728 31358 17740
rect 33965 17731 34023 17737
rect 33965 17728 33977 17731
rect 31352 17700 33977 17728
rect 31352 17688 31358 17700
rect 33965 17697 33977 17700
rect 34011 17728 34023 17731
rect 37826 17728 37832 17740
rect 34011 17700 37832 17728
rect 34011 17697 34023 17700
rect 33965 17691 34023 17697
rect 37826 17688 37832 17700
rect 37884 17688 37890 17740
rect 26878 17620 26884 17672
rect 26936 17660 26942 17672
rect 33689 17663 33747 17669
rect 33689 17660 33701 17663
rect 26936 17632 33701 17660
rect 26936 17620 26942 17632
rect 33689 17629 33701 17632
rect 33735 17629 33747 17663
rect 33689 17623 33747 17629
rect 33778 17484 33784 17536
rect 33836 17524 33842 17536
rect 33836 17496 33881 17524
rect 33836 17484 33842 17496
rect 1104 17434 118864 17456
rect 1104 17382 30398 17434
rect 30450 17382 30462 17434
rect 30514 17382 30526 17434
rect 30578 17382 30590 17434
rect 30642 17382 30654 17434
rect 30706 17382 59846 17434
rect 59898 17382 59910 17434
rect 59962 17382 59974 17434
rect 60026 17382 60038 17434
rect 60090 17382 60102 17434
rect 60154 17382 89294 17434
rect 89346 17382 89358 17434
rect 89410 17382 89422 17434
rect 89474 17382 89486 17434
rect 89538 17382 89550 17434
rect 89602 17382 118864 17434
rect 1104 17360 118864 17382
rect 59722 17280 59728 17332
rect 59780 17320 59786 17332
rect 70118 17320 70124 17332
rect 59780 17292 70124 17320
rect 59780 17280 59786 17292
rect 70118 17280 70124 17292
rect 70176 17280 70182 17332
rect 65978 17212 65984 17264
rect 66036 17252 66042 17264
rect 115198 17252 115204 17264
rect 66036 17224 115204 17252
rect 66036 17212 66042 17224
rect 115198 17212 115204 17224
rect 115256 17212 115262 17264
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 1946 17184 1952 17196
rect 1627 17156 1952 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 82906 17184 82912 17196
rect 82867 17156 82912 17184
rect 82906 17144 82912 17156
rect 82964 17144 82970 17196
rect 1394 17048 1400 17060
rect 1355 17020 1400 17048
rect 1394 17008 1400 17020
rect 1452 17008 1458 17060
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 82725 16983 82783 16989
rect 82725 16949 82737 16983
rect 82771 16980 82783 16983
rect 90358 16980 90364 16992
rect 82771 16952 90364 16980
rect 82771 16949 82783 16952
rect 82725 16943 82783 16949
rect 90358 16940 90364 16952
rect 90416 16940 90422 16992
rect 1104 16890 118864 16912
rect 1104 16838 15674 16890
rect 15726 16838 15738 16890
rect 15790 16838 15802 16890
rect 15854 16838 15866 16890
rect 15918 16838 15930 16890
rect 15982 16838 45122 16890
rect 45174 16838 45186 16890
rect 45238 16838 45250 16890
rect 45302 16838 45314 16890
rect 45366 16838 45378 16890
rect 45430 16838 74570 16890
rect 74622 16838 74634 16890
rect 74686 16838 74698 16890
rect 74750 16838 74762 16890
rect 74814 16838 74826 16890
rect 74878 16838 104018 16890
rect 104070 16838 104082 16890
rect 104134 16838 104146 16890
rect 104198 16838 104210 16890
rect 104262 16838 104274 16890
rect 104326 16838 118864 16890
rect 1104 16816 118864 16838
rect 25406 16668 25412 16720
rect 25464 16708 25470 16720
rect 81805 16711 81863 16717
rect 81805 16708 81817 16711
rect 25464 16680 81817 16708
rect 25464 16668 25470 16680
rect 81805 16677 81817 16680
rect 81851 16708 81863 16711
rect 81851 16680 82492 16708
rect 81851 16677 81863 16680
rect 81805 16671 81863 16677
rect 3510 16600 3516 16652
rect 3568 16640 3574 16652
rect 71501 16643 71559 16649
rect 71501 16640 71513 16643
rect 3568 16612 71513 16640
rect 3568 16600 3574 16612
rect 71501 16609 71513 16612
rect 71547 16609 71559 16643
rect 71501 16603 71559 16609
rect 1578 16572 1584 16584
rect 1539 16544 1584 16572
rect 1578 16532 1584 16544
rect 1636 16532 1642 16584
rect 66901 16575 66959 16581
rect 66901 16541 66913 16575
rect 66947 16572 66959 16575
rect 70578 16572 70584 16584
rect 66947 16544 70584 16572
rect 66947 16541 66959 16544
rect 66901 16535 66959 16541
rect 70578 16532 70584 16544
rect 70636 16532 70642 16584
rect 82464 16572 82492 16680
rect 83292 16680 103514 16708
rect 82722 16640 82728 16652
rect 82683 16612 82728 16640
rect 82722 16600 82728 16612
rect 82780 16600 82786 16652
rect 83292 16649 83320 16680
rect 83277 16643 83335 16649
rect 83277 16640 83289 16643
rect 83187 16612 83289 16640
rect 83277 16609 83289 16612
rect 83323 16609 83335 16643
rect 103486 16640 103514 16680
rect 117593 16643 117651 16649
rect 117593 16640 117605 16643
rect 103486 16612 117605 16640
rect 83277 16603 83335 16609
rect 117593 16609 117605 16612
rect 117639 16609 117651 16643
rect 117593 16603 117651 16609
rect 82633 16575 82691 16581
rect 82633 16572 82645 16575
rect 82464 16544 82645 16572
rect 82633 16541 82645 16544
rect 82679 16541 82691 16575
rect 82633 16535 82691 16541
rect 2590 16504 2596 16516
rect 1412 16476 2596 16504
rect 1412 16445 1440 16476
rect 2590 16464 2596 16476
rect 2648 16464 2654 16516
rect 70762 16464 70768 16516
rect 70820 16504 70826 16516
rect 71225 16507 71283 16513
rect 71225 16504 71237 16507
rect 70820 16476 71237 16504
rect 70820 16464 70826 16476
rect 71225 16473 71237 16476
rect 71271 16473 71283 16507
rect 71225 16467 71283 16473
rect 82541 16507 82599 16513
rect 82541 16473 82553 16507
rect 82587 16504 82599 16507
rect 83292 16504 83320 16603
rect 117222 16532 117228 16584
rect 117280 16572 117286 16584
rect 117317 16575 117375 16581
rect 117317 16572 117329 16575
rect 117280 16544 117329 16572
rect 117280 16532 117286 16544
rect 117317 16541 117329 16544
rect 117363 16541 117375 16575
rect 117317 16535 117375 16541
rect 82587 16476 83320 16504
rect 82587 16473 82599 16476
rect 82541 16467 82599 16473
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16405 1455 16439
rect 1397 16399 1455 16405
rect 1946 16396 1952 16448
rect 2004 16436 2010 16448
rect 67085 16439 67143 16445
rect 67085 16436 67097 16439
rect 2004 16408 67097 16436
rect 2004 16396 2010 16408
rect 67085 16405 67097 16408
rect 67131 16405 67143 16439
rect 67085 16399 67143 16405
rect 82173 16439 82231 16445
rect 82173 16405 82185 16439
rect 82219 16436 82231 16439
rect 82906 16436 82912 16448
rect 82219 16408 82912 16436
rect 82219 16405 82231 16408
rect 82173 16399 82231 16405
rect 82906 16396 82912 16408
rect 82964 16396 82970 16448
rect 1104 16346 118864 16368
rect 1104 16294 30398 16346
rect 30450 16294 30462 16346
rect 30514 16294 30526 16346
rect 30578 16294 30590 16346
rect 30642 16294 30654 16346
rect 30706 16294 59846 16346
rect 59898 16294 59910 16346
rect 59962 16294 59974 16346
rect 60026 16294 60038 16346
rect 60090 16294 60102 16346
rect 60154 16294 89294 16346
rect 89346 16294 89358 16346
rect 89410 16294 89422 16346
rect 89474 16294 89486 16346
rect 89538 16294 89550 16346
rect 89602 16294 118864 16346
rect 1104 16272 118864 16294
rect 68189 16167 68247 16173
rect 68189 16133 68201 16167
rect 68235 16164 68247 16167
rect 68278 16164 68284 16176
rect 68235 16136 68284 16164
rect 68235 16133 68247 16136
rect 68189 16127 68247 16133
rect 68278 16124 68284 16136
rect 68336 16124 68342 16176
rect 66993 16099 67051 16105
rect 66993 16065 67005 16099
rect 67039 16096 67051 16099
rect 67450 16096 67456 16108
rect 67039 16068 67456 16096
rect 67039 16065 67051 16068
rect 66993 16059 67051 16065
rect 67450 16056 67456 16068
rect 67508 16056 67514 16108
rect 68373 16099 68431 16105
rect 68373 16065 68385 16099
rect 68419 16096 68431 16099
rect 68462 16096 68468 16108
rect 68419 16068 68468 16096
rect 68419 16065 68431 16068
rect 68373 16059 68431 16065
rect 68462 16056 68468 16068
rect 68520 16056 68526 16108
rect 69293 16099 69351 16105
rect 69293 16065 69305 16099
rect 69339 16096 69351 16099
rect 69566 16096 69572 16108
rect 69339 16068 69572 16096
rect 69339 16065 69351 16068
rect 69293 16059 69351 16065
rect 69566 16056 69572 16068
rect 69624 16056 69630 16108
rect 66809 15963 66867 15969
rect 66809 15929 66821 15963
rect 66855 15960 66867 15963
rect 68922 15960 68928 15972
rect 66855 15932 68928 15960
rect 66855 15929 66867 15932
rect 66809 15923 66867 15929
rect 68922 15920 68928 15932
rect 68980 15920 68986 15972
rect 68370 15852 68376 15904
rect 68428 15892 68434 15904
rect 68557 15895 68615 15901
rect 68557 15892 68569 15895
rect 68428 15864 68569 15892
rect 68428 15852 68434 15864
rect 68557 15861 68569 15864
rect 68603 15861 68615 15895
rect 68557 15855 68615 15861
rect 69477 15895 69535 15901
rect 69477 15861 69489 15895
rect 69523 15892 69535 15895
rect 70578 15892 70584 15904
rect 69523 15864 70584 15892
rect 69523 15861 69535 15864
rect 69477 15855 69535 15861
rect 70578 15852 70584 15864
rect 70636 15852 70642 15904
rect 118142 15892 118148 15904
rect 118103 15864 118148 15892
rect 118142 15852 118148 15864
rect 118200 15852 118206 15904
rect 1104 15802 118864 15824
rect 1104 15750 15674 15802
rect 15726 15750 15738 15802
rect 15790 15750 15802 15802
rect 15854 15750 15866 15802
rect 15918 15750 15930 15802
rect 15982 15750 45122 15802
rect 45174 15750 45186 15802
rect 45238 15750 45250 15802
rect 45302 15750 45314 15802
rect 45366 15750 45378 15802
rect 45430 15750 74570 15802
rect 74622 15750 74634 15802
rect 74686 15750 74698 15802
rect 74750 15750 74762 15802
rect 74814 15750 74826 15802
rect 74878 15750 104018 15802
rect 104070 15750 104082 15802
rect 104134 15750 104146 15802
rect 104198 15750 104210 15802
rect 104262 15750 104274 15802
rect 104326 15750 118864 15802
rect 1104 15728 118864 15750
rect 68830 15688 68836 15700
rect 67468 15660 68836 15688
rect 53834 15512 53840 15564
rect 53892 15552 53898 15564
rect 66165 15555 66223 15561
rect 66165 15552 66177 15555
rect 53892 15524 66177 15552
rect 53892 15512 53898 15524
rect 66165 15521 66177 15524
rect 66211 15521 66223 15555
rect 66165 15515 66223 15521
rect 67082 15512 67088 15564
rect 67140 15552 67146 15564
rect 67468 15561 67496 15660
rect 68830 15648 68836 15660
rect 68888 15648 68894 15700
rect 69566 15688 69572 15700
rect 69527 15660 69572 15688
rect 69566 15648 69572 15660
rect 69624 15648 69630 15700
rect 70762 15688 70768 15700
rect 70723 15660 70768 15688
rect 70762 15648 70768 15660
rect 70820 15648 70826 15700
rect 67269 15555 67327 15561
rect 67269 15552 67281 15555
rect 67140 15524 67281 15552
rect 67140 15512 67146 15524
rect 67269 15521 67281 15524
rect 67315 15521 67327 15555
rect 67269 15515 67327 15521
rect 67453 15555 67511 15561
rect 67453 15521 67465 15555
rect 67499 15521 67511 15555
rect 67453 15515 67511 15521
rect 68278 15512 68284 15564
rect 68336 15552 68342 15564
rect 71314 15552 71320 15564
rect 68336 15524 68381 15552
rect 71275 15524 71320 15552
rect 68336 15512 68342 15524
rect 71314 15512 71320 15524
rect 71372 15512 71378 15564
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15484 1639 15487
rect 10410 15484 10416 15496
rect 1627 15456 10416 15484
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 56686 15484 56692 15496
rect 45526 15456 56692 15484
rect 30653 15419 30711 15425
rect 30653 15416 30665 15419
rect 26206 15388 30665 15416
rect 1394 15348 1400 15360
rect 1355 15320 1400 15348
rect 1394 15308 1400 15320
rect 1452 15308 1458 15360
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 26206 15348 26234 15388
rect 30653 15385 30665 15388
rect 30699 15385 30711 15419
rect 30653 15379 30711 15385
rect 30837 15419 30895 15425
rect 30837 15385 30849 15419
rect 30883 15416 30895 15419
rect 45526 15416 45554 15456
rect 56686 15444 56692 15456
rect 56744 15444 56750 15496
rect 64877 15487 64935 15493
rect 64877 15453 64889 15487
rect 64923 15484 64935 15487
rect 64966 15484 64972 15496
rect 64923 15456 64972 15484
rect 64923 15453 64935 15456
rect 64877 15447 64935 15453
rect 64966 15444 64972 15456
rect 65024 15444 65030 15496
rect 65978 15484 65984 15496
rect 65939 15456 65984 15484
rect 65978 15444 65984 15456
rect 66036 15444 66042 15496
rect 67174 15484 67180 15496
rect 67135 15456 67180 15484
rect 67174 15444 67180 15456
rect 67232 15444 67238 15496
rect 67361 15487 67419 15493
rect 67361 15453 67373 15487
rect 67407 15484 67419 15487
rect 67726 15484 67732 15496
rect 67407 15456 67732 15484
rect 67407 15453 67419 15456
rect 67361 15447 67419 15453
rect 67726 15444 67732 15456
rect 67784 15444 67790 15496
rect 68186 15484 68192 15496
rect 68147 15456 68192 15484
rect 68186 15444 68192 15456
rect 68244 15444 68250 15496
rect 68373 15487 68431 15493
rect 68373 15453 68385 15487
rect 68419 15453 68431 15487
rect 68373 15447 68431 15453
rect 68465 15487 68523 15493
rect 68465 15453 68477 15487
rect 68511 15453 68523 15487
rect 68465 15447 68523 15453
rect 68925 15487 68983 15493
rect 68925 15453 68937 15487
rect 68971 15484 68983 15487
rect 69198 15484 69204 15496
rect 68971 15456 69204 15484
rect 68971 15453 68983 15456
rect 68925 15447 68983 15453
rect 66073 15419 66131 15425
rect 66073 15416 66085 15419
rect 30883 15388 45554 15416
rect 56152 15388 66085 15416
rect 30883 15385 30895 15388
rect 30837 15379 30895 15385
rect 10928 15320 26234 15348
rect 10928 15308 10934 15320
rect 32766 15308 32772 15360
rect 32824 15348 32830 15360
rect 56152 15348 56180 15388
rect 66073 15385 66085 15388
rect 66119 15416 66131 15419
rect 66625 15419 66683 15425
rect 66625 15416 66637 15419
rect 66119 15388 66637 15416
rect 66119 15385 66131 15388
rect 66073 15379 66131 15385
rect 66625 15385 66637 15388
rect 66671 15385 66683 15419
rect 67744 15416 67772 15444
rect 68388 15416 68416 15447
rect 67744 15388 68416 15416
rect 66625 15379 66683 15385
rect 64690 15348 64696 15360
rect 32824 15320 56180 15348
rect 64651 15320 64696 15348
rect 32824 15308 32830 15320
rect 64690 15308 64696 15320
rect 64748 15308 64754 15360
rect 65613 15351 65671 15357
rect 65613 15317 65625 15351
rect 65659 15348 65671 15351
rect 65794 15348 65800 15360
rect 65659 15320 65800 15348
rect 65659 15317 65671 15320
rect 65613 15311 65671 15317
rect 65794 15308 65800 15320
rect 65852 15308 65858 15360
rect 66990 15348 66996 15360
rect 66951 15320 66996 15348
rect 66990 15308 66996 15320
rect 67048 15308 67054 15360
rect 67542 15308 67548 15360
rect 67600 15348 67606 15360
rect 68005 15351 68063 15357
rect 68005 15348 68017 15351
rect 67600 15320 68017 15348
rect 67600 15308 67606 15320
rect 68005 15317 68017 15320
rect 68051 15317 68063 15351
rect 68480 15348 68508 15447
rect 69198 15444 69204 15456
rect 69256 15484 69262 15496
rect 69256 15456 74534 15484
rect 69256 15444 69262 15456
rect 68738 15376 68744 15428
rect 68796 15416 68802 15428
rect 69385 15419 69443 15425
rect 69385 15416 69397 15419
rect 68796 15388 69397 15416
rect 68796 15376 68802 15388
rect 69385 15385 69397 15388
rect 69431 15416 69443 15419
rect 69658 15416 69664 15428
rect 69431 15388 69664 15416
rect 69431 15385 69443 15388
rect 69385 15379 69443 15385
rect 69658 15376 69664 15388
rect 69716 15376 69722 15428
rect 74506 15416 74534 15456
rect 117406 15416 117412 15428
rect 74506 15388 117412 15416
rect 117406 15376 117412 15388
rect 117464 15376 117470 15428
rect 69750 15348 69756 15360
rect 68480 15320 69756 15348
rect 68005 15311 68063 15317
rect 69750 15308 69756 15320
rect 69808 15308 69814 15360
rect 71130 15348 71136 15360
rect 71091 15320 71136 15348
rect 71130 15308 71136 15320
rect 71188 15308 71194 15360
rect 71225 15351 71283 15357
rect 71225 15317 71237 15351
rect 71271 15348 71283 15351
rect 71869 15351 71927 15357
rect 71869 15348 71881 15351
rect 71271 15320 71881 15348
rect 71271 15317 71283 15320
rect 71225 15311 71283 15317
rect 71869 15317 71881 15320
rect 71915 15348 71927 15351
rect 112530 15348 112536 15360
rect 71915 15320 112536 15348
rect 71915 15317 71927 15320
rect 71869 15311 71927 15317
rect 112530 15308 112536 15320
rect 112588 15308 112594 15360
rect 1104 15258 118864 15280
rect 1104 15206 30398 15258
rect 30450 15206 30462 15258
rect 30514 15206 30526 15258
rect 30578 15206 30590 15258
rect 30642 15206 30654 15258
rect 30706 15206 59846 15258
rect 59898 15206 59910 15258
rect 59962 15206 59974 15258
rect 60026 15206 60038 15258
rect 60090 15206 60102 15258
rect 60154 15206 89294 15258
rect 89346 15206 89358 15258
rect 89410 15206 89422 15258
rect 89474 15206 89486 15258
rect 89538 15206 89550 15258
rect 89602 15206 118864 15258
rect 1104 15184 118864 15206
rect 10410 15104 10416 15156
rect 10468 15144 10474 15156
rect 10505 15147 10563 15153
rect 10505 15144 10517 15147
rect 10468 15116 10517 15144
rect 10468 15104 10474 15116
rect 10505 15113 10517 15116
rect 10551 15113 10563 15147
rect 10505 15107 10563 15113
rect 64874 15104 64880 15156
rect 64932 15144 64938 15156
rect 118050 15144 118056 15156
rect 64932 15116 118056 15144
rect 64932 15104 64938 15116
rect 118050 15104 118056 15116
rect 118108 15104 118114 15156
rect 64138 15036 64144 15088
rect 64196 15076 64202 15088
rect 64233 15079 64291 15085
rect 64233 15076 64245 15079
rect 64196 15048 64245 15076
rect 64196 15036 64202 15048
rect 64233 15045 64245 15048
rect 64279 15045 64291 15079
rect 64233 15039 64291 15045
rect 65058 15036 65064 15088
rect 65116 15076 65122 15088
rect 65153 15079 65211 15085
rect 65153 15076 65165 15079
rect 65116 15048 65165 15076
rect 65116 15036 65122 15048
rect 65153 15045 65165 15048
rect 65199 15045 65211 15079
rect 66530 15076 66536 15088
rect 66491 15048 66536 15076
rect 65153 15039 65211 15045
rect 66530 15036 66536 15048
rect 66588 15076 66594 15088
rect 67361 15079 67419 15085
rect 67361 15076 67373 15079
rect 66588 15048 67373 15076
rect 66588 15036 66594 15048
rect 67361 15045 67373 15048
rect 67407 15076 67419 15079
rect 68738 15076 68744 15088
rect 67407 15048 68744 15076
rect 67407 15045 67419 15048
rect 67361 15039 67419 15045
rect 68738 15036 68744 15048
rect 68796 15036 68802 15088
rect 68830 15036 68836 15088
rect 68888 15076 68894 15088
rect 69477 15079 69535 15085
rect 69477 15076 69489 15079
rect 68888 15048 69489 15076
rect 68888 15036 68894 15048
rect 69477 15045 69489 15048
rect 69523 15045 69535 15079
rect 69477 15039 69535 15045
rect 69658 15036 69664 15088
rect 69716 15076 69722 15088
rect 69753 15079 69811 15085
rect 69753 15076 69765 15079
rect 69716 15048 69765 15076
rect 69716 15036 69722 15048
rect 69753 15045 69765 15048
rect 69799 15045 69811 15079
rect 69753 15039 69811 15045
rect 70578 15036 70584 15088
rect 70636 15076 70642 15088
rect 71222 15076 71228 15088
rect 70636 15048 71228 15076
rect 70636 15036 70642 15048
rect 2406 14968 2412 15020
rect 2464 15008 2470 15020
rect 8021 15011 8079 15017
rect 8021 15008 8033 15011
rect 2464 14980 8033 15008
rect 2464 14968 2470 14980
rect 8021 14977 8033 14980
rect 8067 14977 8079 15011
rect 8021 14971 8079 14977
rect 10689 15011 10747 15017
rect 10689 14977 10701 15011
rect 10735 15008 10747 15011
rect 10870 15008 10876 15020
rect 10735 14980 10876 15008
rect 10735 14977 10747 14980
rect 10689 14971 10747 14977
rect 10870 14968 10876 14980
rect 10928 14968 10934 15020
rect 49605 15011 49663 15017
rect 49605 14977 49617 15011
rect 49651 15008 49663 15011
rect 50433 15011 50491 15017
rect 50433 15008 50445 15011
rect 49651 14980 50445 15008
rect 49651 14977 49663 14980
rect 49605 14971 49663 14977
rect 50433 14977 50445 14980
rect 50479 15008 50491 15011
rect 50522 15008 50528 15020
rect 50479 14980 50528 15008
rect 50479 14977 50491 14980
rect 50433 14971 50491 14977
rect 50522 14968 50528 14980
rect 50580 15008 50586 15020
rect 53745 15011 53803 15017
rect 53745 15008 53757 15011
rect 50580 14980 53757 15008
rect 50580 14968 50586 14980
rect 53745 14977 53757 14980
rect 53791 15008 53803 15011
rect 54849 15011 54907 15017
rect 54849 15008 54861 15011
rect 53791 14980 54861 15008
rect 53791 14977 53803 14980
rect 53745 14971 53803 14977
rect 54849 14977 54861 14980
rect 54895 15008 54907 15011
rect 55861 15011 55919 15017
rect 55861 15008 55873 15011
rect 54895 14980 55873 15008
rect 54895 14977 54907 14980
rect 54849 14971 54907 14977
rect 55861 14977 55873 14980
rect 55907 14977 55919 15011
rect 55861 14971 55919 14977
rect 63957 15011 64015 15017
rect 63957 14977 63969 15011
rect 64003 15008 64015 15011
rect 64690 15008 64696 15020
rect 64003 14980 64696 15008
rect 64003 14977 64015 14980
rect 63957 14971 64015 14977
rect 64690 14968 64696 14980
rect 64748 15008 64754 15020
rect 64877 15011 64935 15017
rect 64877 15008 64889 15011
rect 64748 14980 64889 15008
rect 64748 14968 64754 14980
rect 64877 14977 64889 14980
rect 64923 15008 64935 15011
rect 65886 15008 65892 15020
rect 64923 14980 65892 15008
rect 64923 14977 64935 14980
rect 64877 14971 64935 14977
rect 65886 14968 65892 14980
rect 65944 14968 65950 15020
rect 67269 15011 67327 15017
rect 67269 14977 67281 15011
rect 67315 15008 67327 15011
rect 69198 15008 69204 15020
rect 67315 14980 68968 15008
rect 69159 14980 69204 15008
rect 67315 14977 67327 14980
rect 67269 14971 67327 14977
rect 41322 14900 41328 14952
rect 41380 14940 41386 14952
rect 50617 14943 50675 14949
rect 50617 14940 50629 14943
rect 41380 14912 50629 14940
rect 41380 14900 41386 14912
rect 50617 14909 50629 14912
rect 50663 14909 50675 14943
rect 54570 14940 54576 14952
rect 54531 14912 54576 14940
rect 50617 14903 50675 14909
rect 54570 14900 54576 14912
rect 54628 14900 54634 14952
rect 56134 14940 56140 14952
rect 56095 14912 56140 14940
rect 56134 14900 56140 14912
rect 56192 14900 56198 14952
rect 64138 14900 64144 14952
rect 64196 14940 64202 14952
rect 67545 14943 67603 14949
rect 64196 14912 67036 14940
rect 64196 14900 64202 14912
rect 8205 14875 8263 14881
rect 8205 14841 8217 14875
rect 8251 14872 8263 14875
rect 43346 14872 43352 14884
rect 8251 14844 43352 14872
rect 8251 14841 8263 14844
rect 8205 14835 8263 14841
rect 43346 14832 43352 14844
rect 43404 14832 43410 14884
rect 64966 14832 64972 14884
rect 65024 14872 65030 14884
rect 66901 14875 66959 14881
rect 66901 14872 66913 14875
rect 65024 14844 66913 14872
rect 65024 14832 65030 14844
rect 66901 14841 66913 14844
rect 66947 14841 66959 14875
rect 67008 14872 67036 14912
rect 67545 14909 67557 14943
rect 67591 14940 67603 14943
rect 68462 14940 68468 14952
rect 67591 14912 68468 14940
rect 67591 14909 67603 14912
rect 67545 14903 67603 14909
rect 68462 14900 68468 14912
rect 68520 14900 68526 14952
rect 68646 14872 68652 14884
rect 67008 14844 68652 14872
rect 66901 14835 66959 14841
rect 68646 14832 68652 14844
rect 68704 14832 68710 14884
rect 68741 14875 68799 14881
rect 68741 14841 68753 14875
rect 68787 14872 68799 14875
rect 68830 14872 68836 14884
rect 68787 14844 68836 14872
rect 68787 14841 68799 14844
rect 68741 14835 68799 14841
rect 68830 14832 68836 14844
rect 68888 14832 68894 14884
rect 68940 14872 68968 14980
rect 69198 14968 69204 14980
rect 69256 14968 69262 15020
rect 69290 14968 69296 15020
rect 69348 15008 69354 15020
rect 69937 15011 69995 15017
rect 69348 14980 69393 15008
rect 69348 14968 69354 14980
rect 69937 14977 69949 15011
rect 69983 15008 69995 15011
rect 70394 15008 70400 15020
rect 69983 14980 70400 15008
rect 69983 14977 69995 14980
rect 69937 14971 69995 14977
rect 70394 14968 70400 14980
rect 70452 14968 70458 15020
rect 70780 15017 70808 15048
rect 71222 15036 71228 15048
rect 71280 15036 71286 15088
rect 70765 15011 70823 15017
rect 70765 14977 70777 15011
rect 70811 14977 70823 15011
rect 70765 14971 70823 14977
rect 70949 15011 71007 15017
rect 70949 14977 70961 15011
rect 70995 14977 71007 15011
rect 70949 14971 71007 14977
rect 70026 14940 70032 14952
rect 69216 14912 70032 14940
rect 69216 14872 69244 14912
rect 70026 14900 70032 14912
rect 70084 14900 70090 14952
rect 70964 14940 70992 14971
rect 94958 14940 94964 14952
rect 70136 14912 70992 14940
rect 74506 14912 94964 14940
rect 68940 14844 69244 14872
rect 69290 14832 69296 14884
rect 69348 14872 69354 14884
rect 70136 14872 70164 14912
rect 69348 14844 70164 14872
rect 69348 14832 69354 14844
rect 37826 14764 37832 14816
rect 37884 14804 37890 14816
rect 49697 14807 49755 14813
rect 49697 14804 49709 14807
rect 37884 14776 49709 14804
rect 37884 14764 37890 14776
rect 49697 14773 49709 14776
rect 49743 14773 49755 14807
rect 53834 14804 53840 14816
rect 53795 14776 53840 14804
rect 49697 14767 49755 14773
rect 53834 14764 53840 14776
rect 53892 14764 53898 14816
rect 58526 14764 58532 14816
rect 58584 14804 58590 14816
rect 65978 14804 65984 14816
rect 58584 14776 65984 14804
rect 58584 14764 58590 14776
rect 65978 14764 65984 14776
rect 66036 14764 66042 14816
rect 66070 14764 66076 14816
rect 66128 14804 66134 14816
rect 69014 14804 69020 14816
rect 66128 14776 69020 14804
rect 66128 14764 66134 14776
rect 69014 14764 69020 14776
rect 69072 14804 69078 14816
rect 69842 14804 69848 14816
rect 69072 14776 69848 14804
rect 69072 14764 69078 14776
rect 69842 14764 69848 14776
rect 69900 14764 69906 14816
rect 70136 14813 70164 14844
rect 70210 14832 70216 14884
rect 70268 14872 70274 14884
rect 74506 14872 74534 14912
rect 94958 14900 94964 14912
rect 95016 14900 95022 14952
rect 70268 14844 74534 14872
rect 70268 14832 70274 14844
rect 70121 14807 70179 14813
rect 70121 14773 70133 14807
rect 70167 14773 70179 14807
rect 70302 14804 70308 14816
rect 70263 14776 70308 14804
rect 70121 14767 70179 14773
rect 70302 14764 70308 14776
rect 70360 14764 70366 14816
rect 70578 14764 70584 14816
rect 70636 14804 70642 14816
rect 70857 14807 70915 14813
rect 70857 14804 70869 14807
rect 70636 14776 70869 14804
rect 70636 14764 70642 14776
rect 70857 14773 70869 14776
rect 70903 14773 70915 14807
rect 70857 14767 70915 14773
rect 1104 14714 118864 14736
rect 1104 14662 15674 14714
rect 15726 14662 15738 14714
rect 15790 14662 15802 14714
rect 15854 14662 15866 14714
rect 15918 14662 15930 14714
rect 15982 14662 45122 14714
rect 45174 14662 45186 14714
rect 45238 14662 45250 14714
rect 45302 14662 45314 14714
rect 45366 14662 45378 14714
rect 45430 14662 74570 14714
rect 74622 14662 74634 14714
rect 74686 14662 74698 14714
rect 74750 14662 74762 14714
rect 74814 14662 74826 14714
rect 74878 14662 104018 14714
rect 104070 14662 104082 14714
rect 104134 14662 104146 14714
rect 104198 14662 104210 14714
rect 104262 14662 104274 14714
rect 104326 14662 118864 14714
rect 1104 14640 118864 14662
rect 55490 14600 55496 14612
rect 55451 14572 55496 14600
rect 55490 14560 55496 14572
rect 55548 14560 55554 14612
rect 67082 14560 67088 14612
rect 67140 14600 67146 14612
rect 71593 14603 71651 14609
rect 71593 14600 71605 14603
rect 67140 14572 68140 14600
rect 67140 14560 67146 14572
rect 2225 14535 2283 14541
rect 2225 14501 2237 14535
rect 2271 14501 2283 14535
rect 68112 14532 68140 14572
rect 68572 14572 71605 14600
rect 68572 14532 68600 14572
rect 71593 14569 71605 14572
rect 71639 14569 71651 14603
rect 118050 14600 118056 14612
rect 118011 14572 118056 14600
rect 71593 14563 71651 14569
rect 118050 14560 118056 14572
rect 118108 14560 118114 14612
rect 68112 14504 68600 14532
rect 2225 14495 2283 14501
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 2240 14396 2268 14495
rect 69842 14492 69848 14544
rect 69900 14532 69906 14544
rect 71406 14532 71412 14544
rect 69900 14504 71412 14532
rect 69900 14492 69906 14504
rect 71406 14492 71412 14504
rect 71464 14492 71470 14544
rect 50430 14424 50436 14476
rect 50488 14464 50494 14476
rect 66257 14467 66315 14473
rect 66257 14464 66269 14467
rect 50488 14436 66269 14464
rect 50488 14424 50494 14436
rect 66257 14433 66269 14436
rect 66303 14433 66315 14467
rect 66257 14427 66315 14433
rect 2406 14396 2412 14408
rect 1627 14368 2268 14396
rect 2367 14368 2412 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 50522 14356 50528 14408
rect 50580 14396 50586 14408
rect 50617 14399 50675 14405
rect 50617 14396 50629 14399
rect 50580 14368 50629 14396
rect 50580 14356 50586 14368
rect 50617 14365 50629 14368
rect 50663 14365 50675 14399
rect 50617 14359 50675 14365
rect 54570 14356 54576 14408
rect 54628 14396 54634 14408
rect 55309 14399 55367 14405
rect 55309 14396 55321 14399
rect 54628 14368 55321 14396
rect 54628 14356 54634 14368
rect 55309 14365 55321 14368
rect 55355 14396 55367 14399
rect 64601 14399 64659 14405
rect 55355 14368 58480 14396
rect 55355 14365 55367 14368
rect 55309 14359 55367 14365
rect 1394 14260 1400 14272
rect 1355 14232 1400 14260
rect 1394 14220 1400 14232
rect 1452 14220 1458 14272
rect 50709 14263 50767 14269
rect 50709 14229 50721 14263
rect 50755 14260 50767 14263
rect 50798 14260 50804 14272
rect 50755 14232 50804 14260
rect 50755 14229 50767 14232
rect 50709 14223 50767 14229
rect 50798 14220 50804 14232
rect 50856 14220 50862 14272
rect 58452 14260 58480 14368
rect 64601 14365 64613 14399
rect 64647 14396 64659 14399
rect 65886 14396 65892 14408
rect 64647 14368 65892 14396
rect 64647 14365 64659 14368
rect 64601 14359 64659 14365
rect 65886 14356 65892 14368
rect 65944 14396 65950 14408
rect 65981 14399 66039 14405
rect 65981 14396 65993 14399
rect 65944 14368 65993 14396
rect 65944 14356 65950 14368
rect 65981 14365 65993 14368
rect 66027 14365 66039 14399
rect 65981 14359 66039 14365
rect 64877 14331 64935 14337
rect 64877 14297 64889 14331
rect 64923 14328 64935 14331
rect 66070 14328 66076 14340
rect 64923 14300 66076 14328
rect 64923 14297 64935 14300
rect 64877 14291 64935 14297
rect 66070 14288 66076 14300
rect 66128 14288 66134 14340
rect 64966 14260 64972 14272
rect 58452 14232 64972 14260
rect 64966 14220 64972 14232
rect 65024 14220 65030 14272
rect 66272 14260 66300 14427
rect 69658 14424 69664 14476
rect 69716 14464 69722 14476
rect 70837 14467 70895 14473
rect 70837 14464 70849 14467
rect 69716 14436 70849 14464
rect 69716 14424 69722 14436
rect 70837 14433 70849 14436
rect 70883 14433 70895 14467
rect 70837 14427 70895 14433
rect 66809 14399 66867 14405
rect 66809 14365 66821 14399
rect 66855 14396 66867 14399
rect 68646 14396 68652 14408
rect 66855 14368 68652 14396
rect 66855 14365 66867 14368
rect 66809 14359 66867 14365
rect 68646 14356 68652 14368
rect 68704 14356 68710 14408
rect 71038 14396 71044 14408
rect 68756 14368 70900 14396
rect 70999 14368 71044 14396
rect 67076 14331 67134 14337
rect 67076 14297 67088 14331
rect 67122 14328 67134 14331
rect 67818 14328 67824 14340
rect 67122 14300 67824 14328
rect 67122 14297 67134 14300
rect 67076 14291 67134 14297
rect 67818 14288 67824 14300
rect 67876 14288 67882 14340
rect 68756 14328 68784 14368
rect 68922 14337 68928 14340
rect 68916 14328 68928 14337
rect 68020 14300 68784 14328
rect 68883 14300 68928 14328
rect 68020 14260 68048 14300
rect 68916 14291 68928 14300
rect 68922 14288 68928 14291
rect 68980 14288 68986 14340
rect 69014 14288 69020 14340
rect 69072 14328 69078 14340
rect 70578 14328 70584 14340
rect 69072 14300 70584 14328
rect 69072 14288 69078 14300
rect 70578 14288 70584 14300
rect 70636 14288 70642 14340
rect 70670 14288 70676 14340
rect 70728 14328 70734 14340
rect 70765 14331 70823 14337
rect 70765 14328 70777 14331
rect 70728 14300 70777 14328
rect 70728 14288 70734 14300
rect 70765 14297 70777 14300
rect 70811 14297 70823 14331
rect 70872 14328 70900 14368
rect 71038 14356 71044 14368
rect 71096 14356 71102 14408
rect 71498 14396 71504 14408
rect 71459 14368 71504 14396
rect 71498 14356 71504 14368
rect 71556 14356 71562 14408
rect 117866 14396 117872 14408
rect 117827 14368 117872 14396
rect 117866 14356 117872 14368
rect 117924 14356 117930 14408
rect 90634 14328 90640 14340
rect 70872 14300 90640 14328
rect 70765 14291 70823 14297
rect 90634 14288 90640 14300
rect 90692 14288 90698 14340
rect 66272 14232 68048 14260
rect 68189 14263 68247 14269
rect 68189 14229 68201 14263
rect 68235 14260 68247 14263
rect 68462 14260 68468 14272
rect 68235 14232 68468 14260
rect 68235 14229 68247 14232
rect 68189 14223 68247 14229
rect 68462 14220 68468 14232
rect 68520 14260 68526 14272
rect 69290 14260 69296 14272
rect 68520 14232 69296 14260
rect 68520 14220 68526 14232
rect 69290 14220 69296 14232
rect 69348 14220 69354 14272
rect 70029 14263 70087 14269
rect 70029 14229 70041 14263
rect 70075 14260 70087 14263
rect 70394 14260 70400 14272
rect 70075 14232 70400 14260
rect 70075 14229 70087 14232
rect 70029 14223 70087 14229
rect 70394 14220 70400 14232
rect 70452 14220 70458 14272
rect 70596 14260 70624 14288
rect 70949 14263 71007 14269
rect 70949 14260 70961 14263
rect 70596 14232 70961 14260
rect 70949 14229 70961 14232
rect 70995 14229 71007 14263
rect 70949 14223 71007 14229
rect 1104 14170 118864 14192
rect 1104 14118 30398 14170
rect 30450 14118 30462 14170
rect 30514 14118 30526 14170
rect 30578 14118 30590 14170
rect 30642 14118 30654 14170
rect 30706 14118 59846 14170
rect 59898 14118 59910 14170
rect 59962 14118 59974 14170
rect 60026 14118 60038 14170
rect 60090 14118 60102 14170
rect 60154 14118 89294 14170
rect 89346 14118 89358 14170
rect 89410 14118 89422 14170
rect 89474 14118 89486 14170
rect 89538 14118 89550 14170
rect 89602 14118 118864 14170
rect 1104 14096 118864 14118
rect 56134 14016 56140 14068
rect 56192 14056 56198 14068
rect 65613 14059 65671 14065
rect 56192 14028 60734 14056
rect 56192 14016 56198 14028
rect 60706 13988 60734 14028
rect 65613 14025 65625 14059
rect 65659 14056 65671 14059
rect 65978 14056 65984 14068
rect 65659 14028 65984 14056
rect 65659 14025 65671 14028
rect 65613 14019 65671 14025
rect 65978 14016 65984 14028
rect 66036 14016 66042 14068
rect 67174 14016 67180 14068
rect 67232 14056 67238 14068
rect 69014 14056 69020 14068
rect 67232 14028 69020 14056
rect 67232 14016 67238 14028
rect 69014 14016 69020 14028
rect 69072 14016 69078 14068
rect 71225 14059 71283 14065
rect 71225 14025 71237 14059
rect 71271 14025 71283 14059
rect 71225 14019 71283 14025
rect 66524 13991 66582 13997
rect 60706 13960 66484 13988
rect 65794 13920 65800 13932
rect 65755 13892 65800 13920
rect 65794 13880 65800 13892
rect 65852 13880 65858 13932
rect 66456 13920 66484 13960
rect 66524 13957 66536 13991
rect 66570 13988 66582 13991
rect 69658 13988 69664 14000
rect 66570 13960 69664 13988
rect 66570 13957 66582 13960
rect 66524 13951 66582 13957
rect 69658 13948 69664 13960
rect 69716 13948 69722 14000
rect 69750 13948 69756 14000
rect 69808 13988 69814 14000
rect 71240 13988 71268 14019
rect 71406 14016 71412 14068
rect 71464 14056 71470 14068
rect 85577 14059 85635 14065
rect 85577 14056 85589 14059
rect 71464 14028 85589 14056
rect 71464 14016 71470 14028
rect 85577 14025 85589 14028
rect 85623 14025 85635 14059
rect 86218 14056 86224 14068
rect 86179 14028 86224 14056
rect 85577 14019 85635 14025
rect 69808 13960 71268 13988
rect 85592 13988 85620 14019
rect 86218 14016 86224 14028
rect 86276 14016 86282 14068
rect 118053 14059 118111 14065
rect 118053 14025 118065 14059
rect 118099 14056 118111 14059
rect 118234 14056 118240 14068
rect 118099 14028 118240 14056
rect 118099 14025 118111 14028
rect 118053 14019 118111 14025
rect 118234 14016 118240 14028
rect 118292 14016 118298 14068
rect 86402 13988 86408 14000
rect 85592 13960 86408 13988
rect 69808 13948 69814 13960
rect 86402 13948 86408 13960
rect 86460 13948 86466 14000
rect 68554 13920 68560 13932
rect 66456 13892 68416 13920
rect 68515 13892 68560 13920
rect 66254 13852 66260 13864
rect 66215 13824 66260 13852
rect 66254 13812 66260 13824
rect 66312 13812 66318 13864
rect 68388 13852 68416 13892
rect 68554 13880 68560 13892
rect 68612 13880 68618 13932
rect 68830 13880 68836 13932
rect 68888 13920 68894 13932
rect 70670 13920 70676 13932
rect 68888 13892 70676 13920
rect 68888 13880 68894 13892
rect 70670 13880 70676 13892
rect 70728 13920 70734 13932
rect 71498 13920 71504 13932
rect 70728 13892 71504 13920
rect 70728 13880 70734 13892
rect 71498 13880 71504 13892
rect 71556 13880 71562 13932
rect 107197 13923 107255 13929
rect 84166 13892 93854 13920
rect 69566 13852 69572 13864
rect 68388 13824 69572 13852
rect 69566 13812 69572 13824
rect 69624 13852 69630 13864
rect 69842 13852 69848 13864
rect 69624 13824 69848 13852
rect 69624 13812 69630 13824
rect 69842 13812 69848 13824
rect 69900 13812 69906 13864
rect 70762 13852 70768 13864
rect 70723 13824 70768 13852
rect 70762 13812 70768 13824
rect 70820 13812 70826 13864
rect 81986 13812 81992 13864
rect 82044 13852 82050 13864
rect 84166 13852 84194 13892
rect 86310 13852 86316 13864
rect 82044 13824 84194 13852
rect 86271 13824 86316 13852
rect 82044 13812 82050 13824
rect 86310 13812 86316 13824
rect 86368 13812 86374 13864
rect 86402 13812 86408 13864
rect 86460 13852 86466 13864
rect 93826 13852 93854 13892
rect 107197 13889 107209 13923
rect 107243 13920 107255 13923
rect 108114 13920 108120 13932
rect 107243 13892 108120 13920
rect 107243 13889 107255 13892
rect 107197 13883 107255 13889
rect 108114 13880 108120 13892
rect 108172 13880 108178 13932
rect 117866 13920 117872 13932
rect 117827 13892 117872 13920
rect 117866 13880 117872 13892
rect 117924 13880 117930 13932
rect 107381 13855 107439 13861
rect 107381 13852 107393 13855
rect 86460 13824 86505 13852
rect 93826 13824 107393 13852
rect 86460 13812 86466 13824
rect 107381 13821 107393 13824
rect 107427 13821 107439 13855
rect 107381 13815 107439 13821
rect 48498 13744 48504 13796
rect 48556 13784 48562 13796
rect 57606 13784 57612 13796
rect 48556 13756 57612 13784
rect 48556 13744 48562 13756
rect 57606 13744 57612 13756
rect 57664 13744 57670 13796
rect 70394 13744 70400 13796
rect 70452 13784 70458 13796
rect 71041 13787 71099 13793
rect 71041 13784 71053 13787
rect 70452 13756 71053 13784
rect 70452 13744 70458 13756
rect 71041 13753 71053 13756
rect 71087 13753 71099 13787
rect 71041 13747 71099 13753
rect 67637 13719 67695 13725
rect 67637 13685 67649 13719
rect 67683 13716 67695 13719
rect 68186 13716 68192 13728
rect 67683 13688 68192 13716
rect 67683 13685 67695 13688
rect 67637 13679 67695 13685
rect 68186 13676 68192 13688
rect 68244 13716 68250 13728
rect 68738 13716 68744 13728
rect 68244 13688 68744 13716
rect 68244 13676 68250 13688
rect 68738 13676 68744 13688
rect 68796 13676 68802 13728
rect 69842 13716 69848 13728
rect 69803 13688 69848 13716
rect 69842 13676 69848 13688
rect 69900 13676 69906 13728
rect 85853 13719 85911 13725
rect 85853 13685 85865 13719
rect 85899 13716 85911 13719
rect 86770 13716 86776 13728
rect 85899 13688 86776 13716
rect 85899 13685 85911 13688
rect 85853 13679 85911 13685
rect 86770 13676 86776 13688
rect 86828 13676 86834 13728
rect 1104 13626 118864 13648
rect 1104 13574 15674 13626
rect 15726 13574 15738 13626
rect 15790 13574 15802 13626
rect 15854 13574 15866 13626
rect 15918 13574 15930 13626
rect 15982 13574 45122 13626
rect 45174 13574 45186 13626
rect 45238 13574 45250 13626
rect 45302 13574 45314 13626
rect 45366 13574 45378 13626
rect 45430 13574 74570 13626
rect 74622 13574 74634 13626
rect 74686 13574 74698 13626
rect 74750 13574 74762 13626
rect 74814 13574 74826 13626
rect 74878 13574 104018 13626
rect 104070 13574 104082 13626
rect 104134 13574 104146 13626
rect 104198 13574 104210 13626
rect 104262 13574 104274 13626
rect 104326 13574 118864 13626
rect 1104 13552 118864 13574
rect 68646 13472 68652 13524
rect 68704 13512 68710 13524
rect 68925 13515 68983 13521
rect 68925 13512 68937 13515
rect 68704 13484 68937 13512
rect 68704 13472 68710 13484
rect 68925 13481 68937 13484
rect 68971 13481 68983 13515
rect 68925 13475 68983 13481
rect 70026 13472 70032 13524
rect 70084 13512 70090 13524
rect 70121 13515 70179 13521
rect 70121 13512 70133 13515
rect 70084 13484 70133 13512
rect 70084 13472 70090 13484
rect 70121 13481 70133 13484
rect 70167 13481 70179 13515
rect 70121 13475 70179 13481
rect 67637 13311 67695 13317
rect 67637 13277 67649 13311
rect 67683 13308 67695 13311
rect 69014 13308 69020 13320
rect 67683 13280 69020 13308
rect 67683 13277 67695 13280
rect 67637 13271 67695 13277
rect 69014 13268 69020 13280
rect 69072 13308 69078 13320
rect 69842 13308 69848 13320
rect 69072 13280 69848 13308
rect 69072 13268 69078 13280
rect 69842 13268 69848 13280
rect 69900 13268 69906 13320
rect 70029 13311 70087 13317
rect 70029 13277 70041 13311
rect 70075 13277 70087 13311
rect 86770 13308 86776 13320
rect 86731 13280 86776 13308
rect 70029 13271 70087 13277
rect 1854 13240 1860 13252
rect 1815 13212 1860 13240
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 16022 13200 16028 13252
rect 16080 13240 16086 13252
rect 42978 13240 42984 13252
rect 16080 13212 42984 13240
rect 16080 13200 16086 13212
rect 42978 13200 42984 13212
rect 43036 13200 43042 13252
rect 67726 13200 67732 13252
rect 67784 13240 67790 13252
rect 70044 13240 70072 13271
rect 86770 13268 86776 13280
rect 86828 13268 86834 13320
rect 118142 13308 118148 13320
rect 118103 13280 118148 13308
rect 118142 13268 118148 13280
rect 118200 13268 118206 13320
rect 67784 13212 70072 13240
rect 67784 13200 67790 13212
rect 1949 13175 2007 13181
rect 1949 13141 1961 13175
rect 1995 13172 2007 13175
rect 31110 13172 31116 13184
rect 1995 13144 31116 13172
rect 1995 13141 2007 13144
rect 1949 13135 2007 13141
rect 31110 13132 31116 13144
rect 31168 13132 31174 13184
rect 86586 13172 86592 13184
rect 86547 13144 86592 13172
rect 86586 13132 86592 13144
rect 86644 13132 86650 13184
rect 117958 13172 117964 13184
rect 117919 13144 117964 13172
rect 117958 13132 117964 13144
rect 118016 13132 118022 13184
rect 1104 13082 118864 13104
rect 1104 13030 30398 13082
rect 30450 13030 30462 13082
rect 30514 13030 30526 13082
rect 30578 13030 30590 13082
rect 30642 13030 30654 13082
rect 30706 13030 59846 13082
rect 59898 13030 59910 13082
rect 59962 13030 59974 13082
rect 60026 13030 60038 13082
rect 60090 13030 60102 13082
rect 60154 13030 89294 13082
rect 89346 13030 89358 13082
rect 89410 13030 89422 13082
rect 89474 13030 89486 13082
rect 89538 13030 89550 13082
rect 89602 13030 118864 13082
rect 1104 13008 118864 13030
rect 32122 12968 32128 12980
rect 32083 12940 32128 12968
rect 32122 12928 32128 12940
rect 32180 12928 32186 12980
rect 67637 12971 67695 12977
rect 67637 12937 67649 12971
rect 67683 12968 67695 12971
rect 67726 12968 67732 12980
rect 67683 12940 67732 12968
rect 67683 12937 67695 12940
rect 67637 12931 67695 12937
rect 67726 12928 67732 12940
rect 67784 12928 67790 12980
rect 67818 12928 67824 12980
rect 67876 12968 67882 12980
rect 68189 12971 68247 12977
rect 68189 12968 68201 12971
rect 67876 12940 68201 12968
rect 67876 12928 67882 12940
rect 68189 12937 68201 12940
rect 68235 12937 68247 12971
rect 68189 12931 68247 12937
rect 69937 12971 69995 12977
rect 69937 12937 69949 12971
rect 69983 12968 69995 12971
rect 71038 12968 71044 12980
rect 69983 12940 71044 12968
rect 69983 12937 69995 12940
rect 69937 12931 69995 12937
rect 71038 12928 71044 12940
rect 71096 12928 71102 12980
rect 73798 12928 73804 12980
rect 73856 12968 73862 12980
rect 76745 12971 76803 12977
rect 76745 12968 76757 12971
rect 73856 12940 76757 12968
rect 73856 12928 73862 12940
rect 76745 12937 76757 12940
rect 76791 12937 76803 12971
rect 76745 12931 76803 12937
rect 66524 12903 66582 12909
rect 66524 12869 66536 12903
rect 66570 12900 66582 12903
rect 66990 12900 66996 12912
rect 66570 12872 66996 12900
rect 66570 12869 66582 12872
rect 66524 12863 66582 12869
rect 66990 12860 66996 12872
rect 67048 12860 67054 12912
rect 70302 12900 70308 12912
rect 68480 12872 70308 12900
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 20622 12832 20628 12844
rect 1627 12804 20628 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 32306 12832 32312 12844
rect 32267 12804 32312 12832
rect 32306 12792 32312 12804
rect 32364 12792 32370 12844
rect 66254 12832 66260 12844
rect 66215 12804 66260 12832
rect 66254 12792 66260 12804
rect 66312 12792 66318 12844
rect 68370 12832 68376 12844
rect 68331 12804 68376 12832
rect 68370 12792 68376 12804
rect 68428 12792 68434 12844
rect 68480 12841 68508 12872
rect 70302 12860 70308 12872
rect 70360 12860 70366 12912
rect 68465 12835 68523 12841
rect 68465 12801 68477 12835
rect 68511 12801 68523 12835
rect 68465 12795 68523 12801
rect 68738 12792 68744 12844
rect 68796 12832 68802 12844
rect 69477 12835 69535 12841
rect 69477 12832 69489 12835
rect 68796 12804 69489 12832
rect 68796 12792 68802 12804
rect 69477 12801 69489 12804
rect 69523 12801 69535 12835
rect 69477 12795 69535 12801
rect 108114 12792 108120 12844
rect 108172 12832 108178 12844
rect 108209 12835 108267 12841
rect 108209 12832 108221 12835
rect 108172 12804 108221 12832
rect 108172 12792 108178 12804
rect 108209 12801 108221 12804
rect 108255 12801 108267 12835
rect 108209 12795 108267 12801
rect 67266 12724 67272 12776
rect 67324 12764 67330 12776
rect 68557 12767 68615 12773
rect 68557 12764 68569 12767
rect 67324 12736 68569 12764
rect 67324 12724 67330 12736
rect 68557 12733 68569 12736
rect 68603 12733 68615 12767
rect 68557 12727 68615 12733
rect 68649 12767 68707 12773
rect 68649 12733 68661 12767
rect 68695 12764 68707 12767
rect 68830 12764 68836 12776
rect 68695 12736 68836 12764
rect 68695 12733 68707 12736
rect 68649 12727 68707 12733
rect 68830 12724 68836 12736
rect 68888 12724 68894 12776
rect 76837 12767 76895 12773
rect 76837 12733 76849 12767
rect 76883 12733 76895 12767
rect 77018 12764 77024 12776
rect 76979 12736 77024 12764
rect 76837 12727 76895 12733
rect 76101 12699 76159 12705
rect 76101 12665 76113 12699
rect 76147 12696 76159 12699
rect 76852 12696 76880 12727
rect 77018 12724 77024 12736
rect 77076 12724 77082 12776
rect 76147 12668 76880 12696
rect 76147 12665 76159 12668
rect 76101 12659 76159 12665
rect 1394 12628 1400 12640
rect 1355 12600 1400 12628
rect 1394 12588 1400 12600
rect 1452 12588 1458 12640
rect 68278 12588 68284 12640
rect 68336 12628 68342 12640
rect 69569 12631 69627 12637
rect 69569 12628 69581 12631
rect 68336 12600 69581 12628
rect 68336 12588 68342 12600
rect 69569 12597 69581 12600
rect 69615 12597 69627 12631
rect 76374 12628 76380 12640
rect 76335 12600 76380 12628
rect 69569 12591 69627 12597
rect 76374 12588 76380 12600
rect 76432 12588 76438 12640
rect 76852 12628 76880 12668
rect 99374 12628 99380 12640
rect 76852 12600 99380 12628
rect 99374 12588 99380 12600
rect 99432 12588 99438 12640
rect 108025 12631 108083 12637
rect 108025 12597 108037 12631
rect 108071 12628 108083 12631
rect 118142 12628 118148 12640
rect 108071 12600 118148 12628
rect 108071 12597 108083 12600
rect 108025 12591 108083 12597
rect 118142 12588 118148 12600
rect 118200 12588 118206 12640
rect 1104 12538 118864 12560
rect 1104 12486 15674 12538
rect 15726 12486 15738 12538
rect 15790 12486 15802 12538
rect 15854 12486 15866 12538
rect 15918 12486 15930 12538
rect 15982 12486 45122 12538
rect 45174 12486 45186 12538
rect 45238 12486 45250 12538
rect 45302 12486 45314 12538
rect 45366 12486 45378 12538
rect 45430 12486 74570 12538
rect 74622 12486 74634 12538
rect 74686 12486 74698 12538
rect 74750 12486 74762 12538
rect 74814 12486 74826 12538
rect 74878 12486 104018 12538
rect 104070 12486 104082 12538
rect 104134 12486 104146 12538
rect 104198 12486 104210 12538
rect 104262 12486 104274 12538
rect 104326 12486 118864 12538
rect 1104 12464 118864 12486
rect 20622 12384 20628 12436
rect 20680 12424 20686 12436
rect 21453 12427 21511 12433
rect 21453 12424 21465 12427
rect 20680 12396 21465 12424
rect 20680 12384 20686 12396
rect 21453 12393 21465 12396
rect 21499 12393 21511 12427
rect 21453 12387 21511 12393
rect 31205 12427 31263 12433
rect 31205 12393 31217 12427
rect 31251 12424 31263 12427
rect 32306 12424 32312 12436
rect 31251 12396 32312 12424
rect 31251 12393 31263 12396
rect 31205 12387 31263 12393
rect 32306 12384 32312 12396
rect 32364 12384 32370 12436
rect 67174 12384 67180 12436
rect 67232 12424 67238 12436
rect 67269 12427 67327 12433
rect 67269 12424 67281 12427
rect 67232 12396 67281 12424
rect 67232 12384 67238 12396
rect 67269 12393 67281 12396
rect 67315 12393 67327 12427
rect 67450 12424 67456 12436
rect 67411 12396 67456 12424
rect 67269 12387 67327 12393
rect 67450 12384 67456 12396
rect 67508 12384 67514 12436
rect 68278 12424 68284 12436
rect 68239 12396 68284 12424
rect 68278 12384 68284 12396
rect 68336 12384 68342 12436
rect 39390 12356 39396 12368
rect 22756 12328 39396 12356
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 22756 12297 22784 12328
rect 39390 12316 39396 12328
rect 39448 12356 39454 12368
rect 41322 12356 41328 12368
rect 39448 12328 41328 12356
rect 39448 12316 39454 12328
rect 41322 12316 41328 12328
rect 41380 12316 41386 12368
rect 22557 12291 22615 12297
rect 22557 12288 22569 12291
rect 11756 12260 22569 12288
rect 11756 12248 11762 12260
rect 22557 12257 22569 12260
rect 22603 12257 22615 12291
rect 22557 12251 22615 12257
rect 22741 12291 22799 12297
rect 22741 12257 22753 12291
rect 22787 12257 22799 12291
rect 22741 12251 22799 12257
rect 31849 12291 31907 12297
rect 31849 12257 31861 12291
rect 31895 12288 31907 12291
rect 31895 12260 41414 12288
rect 31895 12257 31907 12260
rect 31849 12251 31907 12257
rect 21637 12223 21695 12229
rect 21637 12189 21649 12223
rect 21683 12220 21695 12223
rect 21683 12192 22140 12220
rect 21683 12189 21695 12192
rect 21637 12183 21695 12189
rect 22112 12093 22140 12192
rect 29730 12180 29736 12232
rect 29788 12220 29794 12232
rect 31573 12223 31631 12229
rect 31573 12220 31585 12223
rect 29788 12192 31585 12220
rect 29788 12180 29794 12192
rect 31573 12189 31585 12192
rect 31619 12189 31631 12223
rect 41386 12220 41414 12260
rect 43717 12223 43775 12229
rect 43717 12220 43729 12223
rect 41386 12192 43729 12220
rect 31573 12183 31631 12189
rect 43717 12189 43729 12192
rect 43763 12220 43775 12223
rect 55490 12220 55496 12232
rect 43763 12192 55496 12220
rect 43763 12189 43775 12192
rect 43717 12183 43775 12189
rect 55490 12180 55496 12192
rect 55548 12180 55554 12232
rect 67821 12223 67879 12229
rect 67821 12189 67833 12223
rect 67867 12220 67879 12223
rect 68189 12223 68247 12229
rect 68189 12220 68201 12223
rect 67867 12192 68201 12220
rect 67867 12189 67879 12192
rect 67821 12183 67879 12189
rect 68189 12189 68201 12192
rect 68235 12220 68247 12223
rect 70762 12220 70768 12232
rect 68235 12192 70768 12220
rect 68235 12189 68247 12192
rect 68189 12183 68247 12189
rect 70762 12180 70768 12192
rect 70820 12220 70826 12232
rect 71682 12220 71688 12232
rect 70820 12192 71688 12220
rect 70820 12180 70826 12192
rect 71682 12180 71688 12192
rect 71740 12180 71746 12232
rect 22465 12155 22523 12161
rect 22465 12121 22477 12155
rect 22511 12152 22523 12155
rect 23290 12152 23296 12164
rect 22511 12124 23296 12152
rect 22511 12121 22523 12124
rect 22465 12115 22523 12121
rect 23290 12112 23296 12124
rect 23348 12112 23354 12164
rect 31665 12155 31723 12161
rect 31665 12152 31677 12155
rect 30852 12124 31677 12152
rect 30852 12096 30880 12124
rect 31665 12121 31677 12124
rect 31711 12121 31723 12155
rect 43990 12152 43996 12164
rect 43951 12124 43996 12152
rect 31665 12115 31723 12121
rect 43990 12112 43996 12124
rect 44048 12112 44054 12164
rect 67082 12152 67088 12164
rect 67043 12124 67088 12152
rect 67082 12112 67088 12124
rect 67140 12112 67146 12164
rect 67301 12155 67359 12161
rect 67301 12121 67313 12155
rect 67347 12152 67359 12155
rect 67542 12152 67548 12164
rect 67347 12124 67548 12152
rect 67347 12121 67359 12124
rect 67301 12115 67359 12121
rect 67542 12112 67548 12124
rect 67600 12112 67606 12164
rect 22097 12087 22155 12093
rect 22097 12053 22109 12087
rect 22143 12053 22155 12087
rect 30834 12084 30840 12096
rect 30795 12056 30840 12084
rect 22097 12047 22155 12053
rect 30834 12044 30840 12056
rect 30892 12044 30898 12096
rect 71406 12044 71412 12096
rect 71464 12084 71470 12096
rect 87230 12084 87236 12096
rect 71464 12056 87236 12084
rect 71464 12044 71470 12056
rect 87230 12044 87236 12056
rect 87288 12044 87294 12096
rect 1104 11994 118864 12016
rect 1104 11942 30398 11994
rect 30450 11942 30462 11994
rect 30514 11942 30526 11994
rect 30578 11942 30590 11994
rect 30642 11942 30654 11994
rect 30706 11942 59846 11994
rect 59898 11942 59910 11994
rect 59962 11942 59974 11994
rect 60026 11942 60038 11994
rect 60090 11942 60102 11994
rect 60154 11942 89294 11994
rect 89346 11942 89358 11994
rect 89410 11942 89422 11994
rect 89474 11942 89486 11994
rect 89538 11942 89550 11994
rect 89602 11942 118864 11994
rect 1104 11920 118864 11942
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 30834 11880 30840 11892
rect 7892 11852 30840 11880
rect 7892 11840 7898 11852
rect 30834 11840 30840 11852
rect 30892 11840 30898 11892
rect 38470 11840 38476 11892
rect 38528 11880 38534 11892
rect 39209 11883 39267 11889
rect 39209 11880 39221 11883
rect 38528 11852 39221 11880
rect 38528 11840 38534 11852
rect 39209 11849 39221 11852
rect 39255 11849 39267 11883
rect 39209 11843 39267 11849
rect 75546 11840 75552 11892
rect 75604 11880 75610 11892
rect 95234 11880 95240 11892
rect 75604 11852 95240 11880
rect 75604 11840 75610 11852
rect 95234 11840 95240 11852
rect 95292 11840 95298 11892
rect 76374 11772 76380 11824
rect 76432 11812 76438 11824
rect 76929 11815 76987 11821
rect 76929 11812 76941 11815
rect 76432 11784 76941 11812
rect 76432 11772 76438 11784
rect 76929 11781 76941 11784
rect 76975 11781 76987 11815
rect 99650 11812 99656 11824
rect 76929 11775 76987 11781
rect 80026 11784 99656 11812
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1544 11716 1593 11744
rect 1544 11704 1550 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 71682 11704 71688 11756
rect 71740 11744 71746 11756
rect 80026 11744 80054 11784
rect 99650 11772 99656 11784
rect 99708 11772 99714 11824
rect 71740 11716 80054 11744
rect 71740 11704 71746 11716
rect 39301 11679 39359 11685
rect 39301 11676 39313 11679
rect 38488 11648 39313 11676
rect 1394 11608 1400 11620
rect 1355 11580 1400 11608
rect 1394 11568 1400 11580
rect 1452 11568 1458 11620
rect 38488 11552 38516 11648
rect 39301 11645 39313 11648
rect 39347 11645 39359 11679
rect 39301 11639 39359 11645
rect 39390 11636 39396 11688
rect 39448 11676 39454 11688
rect 39448 11648 39493 11676
rect 39448 11636 39454 11648
rect 43990 11636 43996 11688
rect 44048 11676 44054 11688
rect 77018 11676 77024 11688
rect 44048 11648 77024 11676
rect 44048 11636 44054 11648
rect 77018 11636 77024 11648
rect 77076 11636 77082 11688
rect 117314 11676 117320 11688
rect 117275 11648 117320 11676
rect 117314 11636 117320 11648
rect 117372 11636 117378 11688
rect 117406 11636 117412 11688
rect 117464 11676 117470 11688
rect 117593 11679 117651 11685
rect 117593 11676 117605 11679
rect 117464 11648 117605 11676
rect 117464 11636 117470 11648
rect 117593 11645 117605 11648
rect 117639 11645 117651 11679
rect 117593 11639 117651 11645
rect 38470 11540 38476 11552
rect 38431 11512 38476 11540
rect 38470 11500 38476 11512
rect 38528 11500 38534 11552
rect 38841 11543 38899 11549
rect 38841 11509 38853 11543
rect 38887 11540 38899 11543
rect 42518 11540 42524 11552
rect 38887 11512 42524 11540
rect 38887 11509 38899 11512
rect 38841 11503 38899 11509
rect 42518 11500 42524 11512
rect 42576 11500 42582 11552
rect 77021 11543 77079 11549
rect 77021 11509 77033 11543
rect 77067 11540 77079 11543
rect 118142 11540 118148 11552
rect 77067 11512 118148 11540
rect 77067 11509 77079 11512
rect 77021 11503 77079 11509
rect 118142 11500 118148 11512
rect 118200 11500 118206 11552
rect 1104 11450 118864 11472
rect 1104 11398 15674 11450
rect 15726 11398 15738 11450
rect 15790 11398 15802 11450
rect 15854 11398 15866 11450
rect 15918 11398 15930 11450
rect 15982 11398 45122 11450
rect 45174 11398 45186 11450
rect 45238 11398 45250 11450
rect 45302 11398 45314 11450
rect 45366 11398 45378 11450
rect 45430 11398 74570 11450
rect 74622 11398 74634 11450
rect 74686 11398 74698 11450
rect 74750 11398 74762 11450
rect 74814 11398 74826 11450
rect 74878 11398 104018 11450
rect 104070 11398 104082 11450
rect 104134 11398 104146 11450
rect 104198 11398 104210 11450
rect 104262 11398 104274 11450
rect 104326 11398 118864 11450
rect 1104 11376 118864 11398
rect 117958 11268 117964 11280
rect 117919 11240 117964 11268
rect 117958 11228 117964 11240
rect 118016 11228 118022 11280
rect 9214 11200 9220 11212
rect 9175 11172 9220 11200
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 42518 11200 42524 11212
rect 42479 11172 42524 11200
rect 42518 11160 42524 11172
rect 42576 11160 42582 11212
rect 2682 11092 2688 11144
rect 2740 11132 2746 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 2740 11104 8953 11132
rect 2740 11092 2746 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 42797 11135 42855 11141
rect 42797 11101 42809 11135
rect 42843 11132 42855 11135
rect 63402 11132 63408 11144
rect 42843 11104 63408 11132
rect 42843 11101 42855 11104
rect 42797 11095 42855 11101
rect 63402 11092 63408 11104
rect 63460 11092 63466 11144
rect 118142 11132 118148 11144
rect 118103 11104 118148 11132
rect 118142 11092 118148 11104
rect 118200 11092 118206 11144
rect 1104 10906 118864 10928
rect 1104 10854 30398 10906
rect 30450 10854 30462 10906
rect 30514 10854 30526 10906
rect 30578 10854 30590 10906
rect 30642 10854 30654 10906
rect 30706 10854 59846 10906
rect 59898 10854 59910 10906
rect 59962 10854 59974 10906
rect 60026 10854 60038 10906
rect 60090 10854 60102 10906
rect 60154 10854 89294 10906
rect 89346 10854 89358 10906
rect 89410 10854 89422 10906
rect 89474 10854 89486 10906
rect 89538 10854 89550 10906
rect 89602 10854 118864 10906
rect 1104 10832 118864 10854
rect 66254 10752 66260 10804
rect 66312 10792 66318 10804
rect 66349 10795 66407 10801
rect 66349 10792 66361 10795
rect 66312 10764 66361 10792
rect 66312 10752 66318 10764
rect 66349 10761 66361 10764
rect 66395 10761 66407 10795
rect 66349 10755 66407 10761
rect 30926 10684 30932 10736
rect 30984 10724 30990 10736
rect 65061 10727 65119 10733
rect 30984 10696 60734 10724
rect 30984 10684 30990 10696
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 2498 10656 2504 10668
rect 1627 10628 2504 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 60706 10656 60734 10696
rect 65061 10693 65073 10727
rect 65107 10724 65119 10727
rect 69014 10724 69020 10736
rect 65107 10696 69020 10724
rect 65107 10693 65119 10696
rect 65061 10687 65119 10693
rect 69014 10684 69020 10696
rect 69072 10684 69078 10736
rect 82538 10724 82544 10736
rect 70366 10696 82544 10724
rect 70366 10656 70394 10696
rect 82538 10684 82544 10696
rect 82596 10684 82602 10736
rect 60706 10628 70394 10656
rect 36538 10548 36544 10600
rect 36596 10588 36602 10600
rect 91922 10588 91928 10600
rect 36596 10560 91928 10588
rect 36596 10548 36602 10560
rect 91922 10548 91928 10560
rect 91980 10548 91986 10600
rect 32950 10480 32956 10532
rect 33008 10520 33014 10532
rect 105538 10520 105544 10532
rect 33008 10492 105544 10520
rect 33008 10480 33014 10492
rect 105538 10480 105544 10492
rect 105596 10480 105602 10532
rect 1394 10452 1400 10464
rect 1355 10424 1400 10452
rect 1394 10412 1400 10424
rect 1452 10412 1458 10464
rect 82998 10412 83004 10464
rect 83056 10452 83062 10464
rect 111702 10452 111708 10464
rect 83056 10424 111708 10452
rect 83056 10412 83062 10424
rect 111702 10412 111708 10424
rect 111760 10412 111766 10464
rect 1104 10362 118864 10384
rect 1104 10310 15674 10362
rect 15726 10310 15738 10362
rect 15790 10310 15802 10362
rect 15854 10310 15866 10362
rect 15918 10310 15930 10362
rect 15982 10310 45122 10362
rect 45174 10310 45186 10362
rect 45238 10310 45250 10362
rect 45302 10310 45314 10362
rect 45366 10310 45378 10362
rect 45430 10310 74570 10362
rect 74622 10310 74634 10362
rect 74686 10310 74698 10362
rect 74750 10310 74762 10362
rect 74814 10310 74826 10362
rect 74878 10310 104018 10362
rect 104070 10310 104082 10362
rect 104134 10310 104146 10362
rect 104198 10310 104210 10362
rect 104262 10310 104274 10362
rect 104326 10310 118864 10362
rect 1104 10288 118864 10310
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 113634 10208 113640 10260
rect 113692 10248 113698 10260
rect 113729 10251 113787 10257
rect 113729 10248 113741 10251
rect 113692 10220 113741 10248
rect 113692 10208 113698 10220
rect 113729 10217 113741 10220
rect 113775 10217 113787 10251
rect 113729 10211 113787 10217
rect 1486 10004 1492 10056
rect 1544 10044 1550 10056
rect 2682 10044 2688 10056
rect 1544 10016 2688 10044
rect 1544 10004 1550 10016
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 115934 10004 115940 10056
rect 115992 10044 115998 10056
rect 118145 10047 118203 10053
rect 118145 10044 118157 10047
rect 115992 10016 118157 10044
rect 115992 10004 115998 10016
rect 118145 10013 118157 10016
rect 118191 10013 118203 10047
rect 118145 10007 118203 10013
rect 1854 9976 1860 9988
rect 1815 9948 1860 9976
rect 1854 9936 1860 9948
rect 1912 9936 1918 9988
rect 2041 9979 2099 9985
rect 2041 9945 2053 9979
rect 2087 9976 2099 9979
rect 113637 9979 113695 9985
rect 2087 9948 6914 9976
rect 2087 9945 2099 9948
rect 2041 9939 2099 9945
rect 6886 9908 6914 9948
rect 113637 9945 113649 9979
rect 113683 9976 113695 9979
rect 114738 9976 114744 9988
rect 113683 9948 114744 9976
rect 113683 9945 113695 9948
rect 113637 9939 113695 9945
rect 114738 9936 114744 9948
rect 114796 9936 114802 9988
rect 31754 9908 31760 9920
rect 6886 9880 31760 9908
rect 31754 9868 31760 9880
rect 31812 9868 31818 9920
rect 117958 9908 117964 9920
rect 117919 9880 117964 9908
rect 117958 9868 117964 9880
rect 118016 9868 118022 9920
rect 1104 9818 118864 9840
rect 1104 9766 30398 9818
rect 30450 9766 30462 9818
rect 30514 9766 30526 9818
rect 30578 9766 30590 9818
rect 30642 9766 30654 9818
rect 30706 9766 59846 9818
rect 59898 9766 59910 9818
rect 59962 9766 59974 9818
rect 60026 9766 60038 9818
rect 60090 9766 60102 9818
rect 60154 9766 89294 9818
rect 89346 9766 89358 9818
rect 89410 9766 89422 9818
rect 89474 9766 89486 9818
rect 89538 9766 89550 9818
rect 89602 9766 118864 9818
rect 1104 9744 118864 9766
rect 68554 9596 68560 9648
rect 68612 9636 68618 9648
rect 115382 9636 115388 9648
rect 68612 9608 115388 9636
rect 68612 9596 68618 9608
rect 115382 9596 115388 9608
rect 115440 9596 115446 9648
rect 114738 9568 114744 9580
rect 114699 9540 114744 9568
rect 114738 9528 114744 9540
rect 114796 9528 114802 9580
rect 114557 9435 114615 9441
rect 114557 9401 114569 9435
rect 114603 9432 114615 9435
rect 115934 9432 115940 9444
rect 114603 9404 115940 9432
rect 114603 9401 114615 9404
rect 114557 9395 114615 9401
rect 115934 9392 115940 9404
rect 115992 9392 115998 9444
rect 1104 9274 118864 9296
rect 1104 9222 15674 9274
rect 15726 9222 15738 9274
rect 15790 9222 15802 9274
rect 15854 9222 15866 9274
rect 15918 9222 15930 9274
rect 15982 9222 45122 9274
rect 45174 9222 45186 9274
rect 45238 9222 45250 9274
rect 45302 9222 45314 9274
rect 45366 9222 45378 9274
rect 45430 9222 74570 9274
rect 74622 9222 74634 9274
rect 74686 9222 74698 9274
rect 74750 9222 74762 9274
rect 74814 9222 74826 9274
rect 74878 9222 104018 9274
rect 104070 9222 104082 9274
rect 104134 9222 104146 9274
rect 104198 9222 104210 9274
rect 104262 9222 104274 9274
rect 104326 9222 118864 9274
rect 1104 9200 118864 9222
rect 76650 8916 76656 8968
rect 76708 8956 76714 8968
rect 113634 8956 113640 8968
rect 76708 8928 113640 8956
rect 76708 8916 76714 8928
rect 113634 8916 113640 8928
rect 113692 8916 113698 8968
rect 1104 8730 118864 8752
rect 1104 8678 30398 8730
rect 30450 8678 30462 8730
rect 30514 8678 30526 8730
rect 30578 8678 30590 8730
rect 30642 8678 30654 8730
rect 30706 8678 59846 8730
rect 59898 8678 59910 8730
rect 59962 8678 59974 8730
rect 60026 8678 60038 8730
rect 60090 8678 60102 8730
rect 60154 8678 89294 8730
rect 89346 8678 89358 8730
rect 89410 8678 89422 8730
rect 89474 8678 89486 8730
rect 89538 8678 89550 8730
rect 89602 8678 118864 8730
rect 1104 8656 118864 8678
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 29733 8483 29791 8489
rect 29733 8480 29745 8483
rect 1627 8452 29745 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 29733 8449 29745 8452
rect 29779 8449 29791 8483
rect 29733 8443 29791 8449
rect 77202 8440 77208 8492
rect 77260 8480 77266 8492
rect 117593 8483 117651 8489
rect 117593 8480 117605 8483
rect 77260 8452 117605 8480
rect 77260 8440 77266 8452
rect 117593 8449 117605 8452
rect 117639 8480 117651 8483
rect 118145 8483 118203 8489
rect 118145 8480 118157 8483
rect 117639 8452 118157 8480
rect 117639 8449 117651 8452
rect 117593 8443 117651 8449
rect 118145 8449 118157 8452
rect 118191 8449 118203 8483
rect 118145 8443 118203 8449
rect 29454 8412 29460 8424
rect 29415 8384 29460 8412
rect 29454 8372 29460 8384
rect 29512 8372 29518 8424
rect 1394 8344 1400 8356
rect 1355 8316 1400 8344
rect 1394 8304 1400 8316
rect 1452 8304 1458 8356
rect 117958 8344 117964 8356
rect 117919 8316 117964 8344
rect 117958 8304 117964 8316
rect 118016 8304 118022 8356
rect 1104 8186 118864 8208
rect 1104 8134 15674 8186
rect 15726 8134 15738 8186
rect 15790 8134 15802 8186
rect 15854 8134 15866 8186
rect 15918 8134 15930 8186
rect 15982 8134 45122 8186
rect 45174 8134 45186 8186
rect 45238 8134 45250 8186
rect 45302 8134 45314 8186
rect 45366 8134 45378 8186
rect 45430 8134 74570 8186
rect 74622 8134 74634 8186
rect 74686 8134 74698 8186
rect 74750 8134 74762 8186
rect 74814 8134 74826 8186
rect 74878 8134 104018 8186
rect 104070 8134 104082 8186
rect 104134 8134 104146 8186
rect 104198 8134 104210 8186
rect 104262 8134 104274 8186
rect 104326 8134 118864 8186
rect 1104 8112 118864 8134
rect 29454 8032 29460 8084
rect 29512 8072 29518 8084
rect 29733 8075 29791 8081
rect 29733 8072 29745 8075
rect 29512 8044 29745 8072
rect 29512 8032 29518 8044
rect 29733 8041 29745 8044
rect 29779 8041 29791 8075
rect 29733 8035 29791 8041
rect 77202 8004 77208 8016
rect 77163 7976 77208 8004
rect 77202 7964 77208 7976
rect 77260 7964 77266 8016
rect 27522 7896 27528 7948
rect 27580 7936 27586 7948
rect 30285 7939 30343 7945
rect 30285 7936 30297 7939
rect 27580 7908 30297 7936
rect 27580 7896 27586 7908
rect 30285 7905 30297 7908
rect 30331 7936 30343 7939
rect 43990 7936 43996 7948
rect 30331 7908 43996 7936
rect 30331 7905 30343 7908
rect 30285 7899 30343 7905
rect 43990 7896 43996 7908
rect 44048 7896 44054 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 1719 7840 6914 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 6886 7800 6914 7840
rect 60706 7840 80054 7868
rect 30101 7803 30159 7809
rect 30101 7800 30113 7803
rect 6886 7772 30113 7800
rect 30101 7769 30113 7772
rect 30147 7769 30159 7803
rect 30101 7763 30159 7769
rect 46934 7760 46940 7812
rect 46992 7800 46998 7812
rect 60706 7800 60734 7840
rect 46992 7772 60734 7800
rect 46992 7760 46998 7772
rect 76466 7760 76472 7812
rect 76524 7800 76530 7812
rect 77021 7803 77079 7809
rect 77021 7800 77033 7803
rect 76524 7772 77033 7800
rect 76524 7760 76530 7772
rect 77021 7769 77033 7772
rect 77067 7769 77079 7803
rect 80026 7800 80054 7840
rect 116210 7800 116216 7812
rect 80026 7772 116216 7800
rect 77021 7763 77079 7769
rect 116210 7760 116216 7772
rect 116268 7760 116274 7812
rect 30193 7735 30251 7741
rect 30193 7701 30205 7735
rect 30239 7732 30251 7735
rect 30837 7735 30895 7741
rect 30837 7732 30849 7735
rect 30239 7704 30849 7732
rect 30239 7701 30251 7704
rect 30193 7695 30251 7701
rect 30837 7701 30849 7704
rect 30883 7732 30895 7735
rect 48314 7732 48320 7744
rect 30883 7704 48320 7732
rect 30883 7701 30895 7704
rect 30837 7695 30895 7701
rect 48314 7692 48320 7704
rect 48372 7692 48378 7744
rect 1104 7642 118864 7664
rect 1104 7590 30398 7642
rect 30450 7590 30462 7642
rect 30514 7590 30526 7642
rect 30578 7590 30590 7642
rect 30642 7590 30654 7642
rect 30706 7590 59846 7642
rect 59898 7590 59910 7642
rect 59962 7590 59974 7642
rect 60026 7590 60038 7642
rect 60090 7590 60102 7642
rect 60154 7590 89294 7642
rect 89346 7590 89358 7642
rect 89410 7590 89422 7642
rect 89474 7590 89486 7642
rect 89538 7590 89550 7642
rect 89602 7590 118864 7642
rect 1104 7568 118864 7590
rect 70486 7488 70492 7540
rect 70544 7528 70550 7540
rect 71314 7528 71320 7540
rect 70544 7500 71320 7528
rect 70544 7488 70550 7500
rect 71314 7488 71320 7500
rect 71372 7488 71378 7540
rect 86221 7395 86279 7401
rect 86221 7361 86233 7395
rect 86267 7392 86279 7395
rect 86954 7392 86960 7404
rect 86267 7364 86960 7392
rect 86267 7361 86279 7364
rect 86221 7355 86279 7361
rect 86954 7352 86960 7364
rect 87012 7352 87018 7404
rect 117958 7392 117964 7404
rect 117919 7364 117964 7392
rect 117958 7352 117964 7364
rect 118016 7352 118022 7404
rect 4798 7148 4804 7200
rect 4856 7188 4862 7200
rect 86313 7191 86371 7197
rect 86313 7188 86325 7191
rect 4856 7160 86325 7188
rect 4856 7148 4862 7160
rect 86313 7157 86325 7160
rect 86359 7157 86371 7191
rect 86313 7151 86371 7157
rect 86954 7148 86960 7200
rect 87012 7188 87018 7200
rect 118053 7191 118111 7197
rect 118053 7188 118065 7191
rect 87012 7160 118065 7188
rect 87012 7148 87018 7160
rect 118053 7157 118065 7160
rect 118099 7157 118111 7191
rect 118053 7151 118111 7157
rect 1104 7098 118864 7120
rect 1104 7046 15674 7098
rect 15726 7046 15738 7098
rect 15790 7046 15802 7098
rect 15854 7046 15866 7098
rect 15918 7046 15930 7098
rect 15982 7046 45122 7098
rect 45174 7046 45186 7098
rect 45238 7046 45250 7098
rect 45302 7046 45314 7098
rect 45366 7046 45378 7098
rect 45430 7046 74570 7098
rect 74622 7046 74634 7098
rect 74686 7046 74698 7098
rect 74750 7046 74762 7098
rect 74814 7046 74826 7098
rect 74878 7046 104018 7098
rect 104070 7046 104082 7098
rect 104134 7046 104146 7098
rect 104198 7046 104210 7098
rect 104262 7046 104274 7098
rect 104326 7046 118864 7098
rect 1104 7024 118864 7046
rect 64598 6876 64604 6928
rect 64656 6916 64662 6928
rect 69474 6916 69480 6928
rect 64656 6888 69480 6916
rect 64656 6876 64662 6888
rect 69474 6876 69480 6888
rect 69532 6876 69538 6928
rect 49878 6740 49884 6792
rect 49936 6780 49942 6792
rect 50341 6783 50399 6789
rect 50341 6780 50353 6783
rect 49936 6752 50353 6780
rect 49936 6740 49942 6752
rect 50341 6749 50353 6752
rect 50387 6749 50399 6783
rect 50341 6743 50399 6749
rect 50062 6604 50068 6656
rect 50120 6644 50126 6656
rect 50157 6647 50215 6653
rect 50157 6644 50169 6647
rect 50120 6616 50169 6644
rect 50120 6604 50126 6616
rect 50157 6613 50169 6616
rect 50203 6613 50215 6647
rect 50157 6607 50215 6613
rect 1104 6554 118864 6576
rect 1104 6502 30398 6554
rect 30450 6502 30462 6554
rect 30514 6502 30526 6554
rect 30578 6502 30590 6554
rect 30642 6502 30654 6554
rect 30706 6502 59846 6554
rect 59898 6502 59910 6554
rect 59962 6502 59974 6554
rect 60026 6502 60038 6554
rect 60090 6502 60102 6554
rect 60154 6502 89294 6554
rect 89346 6502 89358 6554
rect 89410 6502 89422 6554
rect 89474 6502 89486 6554
rect 89538 6502 89550 6554
rect 89602 6502 118864 6554
rect 1104 6480 118864 6502
rect 49878 6440 49884 6452
rect 49839 6412 49884 6440
rect 49878 6400 49884 6412
rect 49936 6400 49942 6452
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 1946 6304 1952 6316
rect 1627 6276 1952 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 49694 6264 49700 6316
rect 49752 6304 49758 6316
rect 50249 6307 50307 6313
rect 50249 6304 50261 6307
rect 49752 6276 50261 6304
rect 49752 6264 49758 6276
rect 50249 6273 50261 6276
rect 50295 6273 50307 6307
rect 50249 6267 50307 6273
rect 50341 6307 50399 6313
rect 50341 6273 50353 6307
rect 50387 6304 50399 6307
rect 86954 6304 86960 6316
rect 50387 6276 51074 6304
rect 86915 6276 86960 6304
rect 50387 6273 50399 6276
rect 50341 6267 50399 6273
rect 50430 6196 50436 6248
rect 50488 6236 50494 6248
rect 51046 6236 51074 6276
rect 86954 6264 86960 6276
rect 87012 6264 87018 6316
rect 117866 6304 117872 6316
rect 117827 6276 117872 6304
rect 117866 6264 117872 6276
rect 117924 6264 117930 6316
rect 50488 6208 50533 6236
rect 51046 6208 113174 6236
rect 50488 6196 50494 6208
rect 1394 6168 1400 6180
rect 1355 6140 1400 6168
rect 1394 6128 1400 6140
rect 1452 6128 1458 6180
rect 59262 6128 59268 6180
rect 59320 6168 59326 6180
rect 110046 6168 110052 6180
rect 59320 6140 110052 6168
rect 59320 6128 59326 6140
rect 110046 6128 110052 6140
rect 110104 6128 110110 6180
rect 113146 6168 113174 6208
rect 118053 6171 118111 6177
rect 118053 6168 118065 6171
rect 113146 6140 118065 6168
rect 118053 6137 118065 6140
rect 118099 6137 118111 6171
rect 118053 6131 118111 6137
rect 1946 6100 1952 6112
rect 1907 6072 1952 6100
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 86773 6103 86831 6109
rect 86773 6069 86785 6103
rect 86819 6100 86831 6103
rect 87230 6100 87236 6112
rect 86819 6072 87236 6100
rect 86819 6069 86831 6072
rect 86773 6063 86831 6069
rect 87230 6060 87236 6072
rect 87288 6060 87294 6112
rect 1104 6010 118864 6032
rect 1104 5958 15674 6010
rect 15726 5958 15738 6010
rect 15790 5958 15802 6010
rect 15854 5958 15866 6010
rect 15918 5958 15930 6010
rect 15982 5958 45122 6010
rect 45174 5958 45186 6010
rect 45238 5958 45250 6010
rect 45302 5958 45314 6010
rect 45366 5958 45378 6010
rect 45430 5958 74570 6010
rect 74622 5958 74634 6010
rect 74686 5958 74698 6010
rect 74750 5958 74762 6010
rect 74814 5958 74826 6010
rect 74878 5958 104018 6010
rect 104070 5958 104082 6010
rect 104134 5958 104146 6010
rect 104198 5958 104210 6010
rect 104262 5958 104274 6010
rect 104326 5958 118864 6010
rect 1104 5936 118864 5958
rect 57422 5652 57428 5704
rect 57480 5692 57486 5704
rect 65886 5692 65892 5704
rect 57480 5664 65892 5692
rect 57480 5652 57486 5664
rect 65886 5652 65892 5664
rect 65944 5652 65950 5704
rect 1854 5624 1860 5636
rect 1815 5596 1860 5624
rect 1854 5584 1860 5596
rect 1912 5584 1918 5636
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 46566 5556 46572 5568
rect 1995 5528 46572 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 46566 5516 46572 5528
rect 46624 5516 46630 5568
rect 1104 5466 118864 5488
rect 1104 5414 30398 5466
rect 30450 5414 30462 5466
rect 30514 5414 30526 5466
rect 30578 5414 30590 5466
rect 30642 5414 30654 5466
rect 30706 5414 59846 5466
rect 59898 5414 59910 5466
rect 59962 5414 59974 5466
rect 60026 5414 60038 5466
rect 60090 5414 60102 5466
rect 60154 5414 89294 5466
rect 89346 5414 89358 5466
rect 89410 5414 89422 5466
rect 89474 5414 89486 5466
rect 89538 5414 89550 5466
rect 89602 5414 118864 5466
rect 1104 5392 118864 5414
rect 82998 5284 83004 5296
rect 82959 5256 83004 5284
rect 82998 5244 83004 5256
rect 83056 5244 83062 5296
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5176 1458 5228
rect 82814 5216 82820 5228
rect 82775 5188 82820 5216
rect 82814 5176 82820 5188
rect 82872 5176 82878 5228
rect 115658 5176 115664 5228
rect 115716 5216 115722 5228
rect 118145 5219 118203 5225
rect 118145 5216 118157 5219
rect 115716 5188 118157 5216
rect 115716 5176 115722 5188
rect 118145 5185 118157 5188
rect 118191 5185 118203 5219
rect 118145 5179 118203 5185
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 61010 5012 61016 5024
rect 1627 4984 61016 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 61010 4972 61016 4984
rect 61068 4972 61074 5024
rect 117958 5012 117964 5024
rect 117919 4984 117964 5012
rect 117958 4972 117964 4984
rect 118016 4972 118022 5024
rect 1104 4922 118864 4944
rect 1104 4870 15674 4922
rect 15726 4870 15738 4922
rect 15790 4870 15802 4922
rect 15854 4870 15866 4922
rect 15918 4870 15930 4922
rect 15982 4870 45122 4922
rect 45174 4870 45186 4922
rect 45238 4870 45250 4922
rect 45302 4870 45314 4922
rect 45366 4870 45378 4922
rect 45430 4870 74570 4922
rect 74622 4870 74634 4922
rect 74686 4870 74698 4922
rect 74750 4870 74762 4922
rect 74814 4870 74826 4922
rect 74878 4870 104018 4922
rect 104070 4870 104082 4922
rect 104134 4870 104146 4922
rect 104198 4870 104210 4922
rect 104262 4870 104274 4922
rect 104326 4870 118864 4922
rect 1104 4848 118864 4870
rect 42610 4564 42616 4616
rect 42668 4604 42674 4616
rect 79226 4604 79232 4616
rect 42668 4576 79232 4604
rect 42668 4564 42674 4576
rect 79226 4564 79232 4576
rect 79284 4604 79290 4616
rect 79321 4607 79379 4613
rect 79321 4604 79333 4607
rect 79284 4576 79333 4604
rect 79284 4564 79290 4576
rect 79321 4573 79333 4576
rect 79367 4604 79379 4607
rect 79781 4607 79839 4613
rect 79781 4604 79793 4607
rect 79367 4576 79793 4604
rect 79367 4573 79379 4576
rect 79321 4567 79379 4573
rect 79781 4573 79793 4576
rect 79827 4573 79839 4607
rect 79781 4567 79839 4573
rect 79965 4539 80023 4545
rect 60706 4508 79456 4536
rect 37642 4428 37648 4480
rect 37700 4468 37706 4480
rect 60706 4468 60734 4508
rect 37700 4440 60734 4468
rect 37700 4428 37706 4440
rect 70578 4428 70584 4480
rect 70636 4468 70642 4480
rect 71406 4468 71412 4480
rect 70636 4440 71412 4468
rect 70636 4428 70642 4440
rect 71406 4428 71412 4440
rect 71464 4428 71470 4480
rect 79428 4468 79456 4508
rect 79965 4505 79977 4539
rect 80011 4536 80023 4539
rect 115658 4536 115664 4548
rect 80011 4508 115664 4536
rect 80011 4505 80023 4508
rect 79965 4499 80023 4505
rect 115658 4496 115664 4508
rect 115716 4496 115722 4548
rect 117774 4536 117780 4548
rect 117735 4508 117780 4536
rect 117774 4496 117780 4508
rect 117832 4496 117838 4548
rect 117869 4471 117927 4477
rect 117869 4468 117881 4471
rect 79428 4440 117881 4468
rect 117869 4437 117881 4440
rect 117915 4437 117927 4471
rect 117869 4431 117927 4437
rect 1104 4378 118864 4400
rect 1104 4326 30398 4378
rect 30450 4326 30462 4378
rect 30514 4326 30526 4378
rect 30578 4326 30590 4378
rect 30642 4326 30654 4378
rect 30706 4326 59846 4378
rect 59898 4326 59910 4378
rect 59962 4326 59974 4378
rect 60026 4326 60038 4378
rect 60090 4326 60102 4378
rect 60154 4326 89294 4378
rect 89346 4326 89358 4378
rect 89410 4326 89422 4378
rect 89474 4326 89486 4378
rect 89538 4326 89550 4378
rect 89602 4326 118864 4378
rect 1104 4304 118864 4326
rect 60645 4267 60703 4273
rect 60645 4233 60657 4267
rect 60691 4233 60703 4267
rect 82630 4264 82636 4276
rect 60645 4227 60703 4233
rect 60752 4236 61148 4264
rect 60660 4196 60688 4227
rect 60752 4196 60780 4236
rect 59188 4168 59676 4196
rect 60660 4168 60780 4196
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1452 4100 1593 4128
rect 1452 4088 1458 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 2590 4128 2596 4140
rect 1820 4100 2596 4128
rect 1820 4088 1826 4100
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 35710 4088 35716 4140
rect 35768 4128 35774 4140
rect 59188 4128 59216 4168
rect 59648 4140 59676 4168
rect 35768 4100 59216 4128
rect 35768 4088 35774 4100
rect 59262 4088 59268 4140
rect 59320 4128 59326 4140
rect 59541 4131 59599 4137
rect 59541 4128 59553 4131
rect 59320 4100 59553 4128
rect 59320 4088 59326 4100
rect 59541 4097 59553 4100
rect 59587 4097 59599 4131
rect 59541 4091 59599 4097
rect 59630 4088 59636 4140
rect 59688 4088 59694 4140
rect 59814 4088 59820 4140
rect 59872 4128 59878 4140
rect 61013 4131 61071 4137
rect 61013 4128 61025 4131
rect 59872 4100 61025 4128
rect 59872 4088 59878 4100
rect 61013 4097 61025 4100
rect 61059 4097 61071 4131
rect 61120 4128 61148 4236
rect 72344 4236 72648 4264
rect 82591 4236 82636 4264
rect 61746 4156 61752 4208
rect 61804 4196 61810 4208
rect 61804 4168 62160 4196
rect 61804 4156 61810 4168
rect 62025 4131 62083 4137
rect 62025 4128 62037 4131
rect 61120 4100 62037 4128
rect 61013 4091 61071 4097
rect 62025 4097 62037 4100
rect 62071 4097 62083 4131
rect 62132 4128 62160 4168
rect 72344 4128 72372 4236
rect 62132 4100 72372 4128
rect 72620 4128 72648 4236
rect 82630 4224 82636 4236
rect 82688 4224 82694 4276
rect 73062 4156 73068 4208
rect 73120 4196 73126 4208
rect 82541 4199 82599 4205
rect 73120 4168 75316 4196
rect 73120 4156 73126 4168
rect 75288 4128 75316 4168
rect 82541 4165 82553 4199
rect 82587 4196 82599 4199
rect 85482 4196 85488 4208
rect 82587 4168 85488 4196
rect 82587 4165 82599 4168
rect 82541 4159 82599 4165
rect 85482 4156 85488 4168
rect 85540 4156 85546 4208
rect 117961 4199 118019 4205
rect 117961 4165 117973 4199
rect 118007 4196 118019 4199
rect 119798 4196 119804 4208
rect 118007 4168 119804 4196
rect 118007 4165 118019 4168
rect 117961 4159 118019 4165
rect 119798 4156 119804 4168
rect 119856 4156 119862 4208
rect 77202 4128 77208 4140
rect 72620 4100 75224 4128
rect 75288 4100 77208 4128
rect 62025 4091 62083 4097
rect 1946 4020 1952 4072
rect 2004 4060 2010 4072
rect 57238 4060 57244 4072
rect 2004 4032 57244 4060
rect 2004 4020 2010 4032
rect 57238 4020 57244 4032
rect 57296 4020 57302 4072
rect 57330 4020 57336 4072
rect 57388 4060 57394 4072
rect 60277 4063 60335 4069
rect 60277 4060 60289 4063
rect 57388 4032 60289 4060
rect 57388 4020 57394 4032
rect 60277 4029 60289 4032
rect 60323 4060 60335 4063
rect 61105 4063 61163 4069
rect 61105 4060 61117 4063
rect 60323 4032 61117 4060
rect 60323 4029 60335 4032
rect 60277 4023 60335 4029
rect 61105 4029 61117 4032
rect 61151 4029 61163 4063
rect 61105 4023 61163 4029
rect 61289 4063 61347 4069
rect 61289 4029 61301 4063
rect 61335 4060 61347 4063
rect 65058 4060 65064 4072
rect 61335 4032 65064 4060
rect 61335 4029 61347 4032
rect 61289 4023 61347 4029
rect 65058 4020 65064 4032
rect 65116 4020 65122 4072
rect 72602 4020 72608 4072
rect 72660 4060 72666 4072
rect 75196 4060 75224 4100
rect 77202 4088 77208 4100
rect 77260 4088 77266 4140
rect 79226 4128 79232 4140
rect 79187 4100 79232 4128
rect 79226 4088 79232 4100
rect 79284 4088 79290 4140
rect 107470 4128 107476 4140
rect 82648 4100 107476 4128
rect 82648 4060 82676 4100
rect 107470 4088 107476 4100
rect 107528 4088 107534 4140
rect 116854 4128 116860 4140
rect 116815 4100 116860 4128
rect 116854 4088 116860 4100
rect 116912 4128 116918 4140
rect 117409 4131 117467 4137
rect 117409 4128 117421 4131
rect 116912 4100 117421 4128
rect 116912 4088 116918 4100
rect 117409 4097 117421 4100
rect 117455 4097 117467 4131
rect 117409 4091 117467 4097
rect 72660 4032 74304 4060
rect 75196 4032 82676 4060
rect 72660 4020 72666 4032
rect 1397 3995 1455 4001
rect 1397 3961 1409 3995
rect 1443 3992 1455 3995
rect 1486 3992 1492 4004
rect 1443 3964 1492 3992
rect 1443 3961 1455 3964
rect 1397 3955 1455 3961
rect 1486 3952 1492 3964
rect 1544 3952 1550 4004
rect 2130 3952 2136 4004
rect 2188 3992 2194 4004
rect 74166 3992 74172 4004
rect 2188 3964 57560 3992
rect 2188 3952 2194 3964
rect 31478 3884 31484 3936
rect 31536 3924 31542 3936
rect 57330 3924 57336 3936
rect 31536 3896 57336 3924
rect 31536 3884 31542 3896
rect 57330 3884 57336 3896
rect 57388 3884 57394 3936
rect 57532 3924 57560 3964
rect 57716 3964 74172 3992
rect 57716 3924 57744 3964
rect 74166 3952 74172 3964
rect 74224 3952 74230 4004
rect 59354 3924 59360 3936
rect 57532 3896 57744 3924
rect 59315 3896 59360 3924
rect 59354 3884 59360 3896
rect 59412 3884 59418 3936
rect 59630 3884 59636 3936
rect 59688 3924 59694 3936
rect 61746 3924 61752 3936
rect 59688 3896 61752 3924
rect 59688 3884 59694 3896
rect 61746 3884 61752 3896
rect 61804 3884 61810 3936
rect 61841 3927 61899 3933
rect 61841 3893 61853 3927
rect 61887 3924 61899 3927
rect 73062 3924 73068 3936
rect 61887 3896 73068 3924
rect 61887 3893 61899 3896
rect 61841 3887 61899 3893
rect 73062 3884 73068 3896
rect 73120 3884 73126 3936
rect 73154 3884 73160 3936
rect 73212 3924 73218 3936
rect 73706 3924 73712 3936
rect 73212 3896 73712 3924
rect 73212 3884 73218 3896
rect 73706 3884 73712 3896
rect 73764 3924 73770 3936
rect 74074 3924 74080 3936
rect 73764 3896 74080 3924
rect 73764 3884 73770 3896
rect 74074 3884 74080 3896
rect 74132 3884 74138 3936
rect 74276 3924 74304 4032
rect 82722 4020 82728 4072
rect 82780 4060 82786 4072
rect 82780 4032 82825 4060
rect 82780 4020 82786 4032
rect 74350 3952 74356 4004
rect 74408 3992 74414 4004
rect 82630 3992 82636 4004
rect 74408 3964 82636 3992
rect 74408 3952 74414 3964
rect 82630 3952 82636 3964
rect 82688 3952 82694 4004
rect 77018 3924 77024 3936
rect 74276 3896 77024 3924
rect 77018 3884 77024 3896
rect 77076 3884 77082 3936
rect 79045 3927 79103 3933
rect 79045 3893 79057 3927
rect 79091 3924 79103 3927
rect 79502 3924 79508 3936
rect 79091 3896 79508 3924
rect 79091 3893 79103 3896
rect 79045 3887 79103 3893
rect 79502 3884 79508 3896
rect 79560 3884 79566 3936
rect 82173 3927 82231 3933
rect 82173 3893 82185 3927
rect 82219 3924 82231 3927
rect 82814 3924 82820 3936
rect 82219 3896 82820 3924
rect 82219 3893 82231 3896
rect 82173 3887 82231 3893
rect 82814 3884 82820 3896
rect 82872 3884 82878 3936
rect 117225 3927 117283 3933
rect 117225 3893 117237 3927
rect 117271 3924 117283 3927
rect 117958 3924 117964 3936
rect 117271 3896 117964 3924
rect 117271 3893 117283 3896
rect 117225 3887 117283 3893
rect 117958 3884 117964 3896
rect 118016 3884 118022 3936
rect 118050 3884 118056 3936
rect 118108 3924 118114 3936
rect 118108 3896 118153 3924
rect 118108 3884 118114 3896
rect 1104 3834 118864 3856
rect 1104 3782 15674 3834
rect 15726 3782 15738 3834
rect 15790 3782 15802 3834
rect 15854 3782 15866 3834
rect 15918 3782 15930 3834
rect 15982 3782 45122 3834
rect 45174 3782 45186 3834
rect 45238 3782 45250 3834
rect 45302 3782 45314 3834
rect 45366 3782 45378 3834
rect 45430 3782 74570 3834
rect 74622 3782 74634 3834
rect 74686 3782 74698 3834
rect 74750 3782 74762 3834
rect 74814 3782 74826 3834
rect 74878 3782 104018 3834
rect 104070 3782 104082 3834
rect 104134 3782 104146 3834
rect 104198 3782 104210 3834
rect 104262 3782 104274 3834
rect 104326 3782 118864 3834
rect 1104 3760 118864 3782
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 45646 3720 45652 3732
rect 5500 3692 45652 3720
rect 5500 3680 5506 3692
rect 45646 3680 45652 3692
rect 45704 3680 45710 3732
rect 56962 3720 56968 3732
rect 45756 3692 56968 3720
rect 40126 3652 40132 3664
rect 22066 3624 40132 3652
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 22066 3584 22094 3624
rect 40126 3612 40132 3624
rect 40184 3612 40190 3664
rect 40681 3655 40739 3661
rect 40681 3621 40693 3655
rect 40727 3652 40739 3655
rect 45756 3652 45784 3692
rect 56962 3680 56968 3692
rect 57020 3680 57026 3732
rect 57054 3680 57060 3732
rect 57112 3720 57118 3732
rect 59630 3720 59636 3732
rect 57112 3692 59492 3720
rect 59591 3692 59636 3720
rect 57112 3680 57118 3692
rect 57974 3652 57980 3664
rect 40727 3624 45784 3652
rect 46216 3624 57980 3652
rect 40727 3621 40739 3624
rect 40681 3615 40739 3621
rect 20772 3556 22094 3584
rect 20772 3544 20778 3556
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 46216 3584 46244 3624
rect 57974 3612 57980 3624
rect 58032 3612 58038 3664
rect 59464 3652 59492 3692
rect 59630 3680 59636 3692
rect 59688 3680 59694 3732
rect 72326 3680 72332 3732
rect 72384 3720 72390 3732
rect 117130 3720 117136 3732
rect 72384 3692 117136 3720
rect 72384 3680 72390 3692
rect 117130 3680 117136 3692
rect 117188 3680 117194 3732
rect 117682 3720 117688 3732
rect 117240 3692 117688 3720
rect 59814 3652 59820 3664
rect 59464 3624 59820 3652
rect 59814 3612 59820 3624
rect 59872 3612 59878 3664
rect 61010 3612 61016 3664
rect 61068 3652 61074 3664
rect 72234 3652 72240 3664
rect 61068 3624 72240 3652
rect 61068 3612 61074 3624
rect 72234 3612 72240 3624
rect 72292 3612 72298 3664
rect 73062 3612 73068 3664
rect 73120 3652 73126 3664
rect 73985 3655 74043 3661
rect 73985 3652 73997 3655
rect 73120 3624 73997 3652
rect 73120 3612 73126 3624
rect 73985 3621 73997 3624
rect 74031 3621 74043 3655
rect 73985 3615 74043 3621
rect 74074 3612 74080 3664
rect 74132 3652 74138 3664
rect 117240 3652 117268 3692
rect 117682 3680 117688 3692
rect 117740 3680 117746 3732
rect 74132 3624 117268 3652
rect 118053 3655 118111 3661
rect 74132 3612 74138 3624
rect 118053 3621 118065 3655
rect 118099 3621 118111 3655
rect 118053 3615 118111 3621
rect 33652 3556 46244 3584
rect 33652 3544 33658 3556
rect 46842 3544 46848 3596
rect 46900 3584 46906 3596
rect 57054 3584 57060 3596
rect 46900 3556 57060 3584
rect 46900 3544 46906 3556
rect 57054 3544 57060 3556
rect 57112 3544 57118 3596
rect 57146 3544 57152 3596
rect 57204 3584 57210 3596
rect 58066 3584 58072 3596
rect 57204 3556 58072 3584
rect 57204 3544 57210 3556
rect 58066 3544 58072 3556
rect 58124 3544 58130 3596
rect 61105 3587 61163 3593
rect 61105 3584 61117 3587
rect 58176 3556 61117 3584
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 2222 3516 2228 3528
rect 2183 3488 2228 3516
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 658 3408 664 3460
rect 716 3448 722 3460
rect 2884 3448 2912 3479
rect 32122 3476 32128 3528
rect 32180 3516 32186 3528
rect 32861 3519 32919 3525
rect 32861 3516 32873 3519
rect 32180 3488 32873 3516
rect 32180 3476 32186 3488
rect 32861 3485 32873 3488
rect 32907 3485 32919 3519
rect 32861 3479 32919 3485
rect 33778 3476 33784 3528
rect 33836 3516 33842 3528
rect 40310 3516 40316 3528
rect 33836 3488 40316 3516
rect 33836 3476 33842 3488
rect 40310 3476 40316 3488
rect 40368 3476 40374 3528
rect 40586 3476 40592 3528
rect 40644 3516 40650 3528
rect 40865 3519 40923 3525
rect 40865 3516 40877 3519
rect 40644 3488 40877 3516
rect 40644 3476 40650 3488
rect 40865 3485 40877 3488
rect 40911 3485 40923 3519
rect 40865 3479 40923 3485
rect 41506 3476 41512 3528
rect 41564 3516 41570 3528
rect 42426 3516 42432 3528
rect 41564 3488 42432 3516
rect 41564 3476 41570 3488
rect 42426 3476 42432 3488
rect 42484 3476 42490 3528
rect 42797 3519 42855 3525
rect 42797 3485 42809 3519
rect 42843 3485 42855 3519
rect 42797 3479 42855 3485
rect 716 3420 2912 3448
rect 716 3408 722 3420
rect 34974 3408 34980 3460
rect 35032 3448 35038 3460
rect 40402 3448 40408 3460
rect 35032 3420 40408 3448
rect 35032 3408 35038 3420
rect 40402 3408 40408 3420
rect 40460 3408 40466 3460
rect 42812 3392 42840 3479
rect 45738 3476 45744 3528
rect 45796 3516 45802 3528
rect 46017 3519 46075 3525
rect 46017 3516 46029 3519
rect 45796 3488 46029 3516
rect 45796 3476 45802 3488
rect 46017 3485 46029 3488
rect 46063 3485 46075 3519
rect 46017 3479 46075 3485
rect 47029 3519 47087 3525
rect 47029 3485 47041 3519
rect 47075 3516 47087 3519
rect 47210 3516 47216 3528
rect 47075 3488 47216 3516
rect 47075 3485 47087 3488
rect 47029 3479 47087 3485
rect 47210 3476 47216 3488
rect 47268 3476 47274 3528
rect 47673 3519 47731 3525
rect 47673 3485 47685 3519
rect 47719 3516 47731 3519
rect 47946 3516 47952 3528
rect 47719 3488 47952 3516
rect 47719 3485 47731 3488
rect 47673 3479 47731 3485
rect 47946 3476 47952 3488
rect 48004 3476 48010 3528
rect 48038 3476 48044 3528
rect 48096 3516 48102 3528
rect 50706 3516 50712 3528
rect 48096 3488 50712 3516
rect 48096 3476 48102 3488
rect 50706 3476 50712 3488
rect 50764 3476 50770 3528
rect 50816 3488 51074 3516
rect 47302 3408 47308 3460
rect 47360 3448 47366 3460
rect 50816 3448 50844 3488
rect 47360 3420 50844 3448
rect 51046 3448 51074 3488
rect 52178 3476 52184 3528
rect 52236 3516 52242 3528
rect 52457 3519 52515 3525
rect 52457 3516 52469 3519
rect 52236 3488 52469 3516
rect 52236 3476 52242 3488
rect 52457 3485 52469 3488
rect 52503 3485 52515 3519
rect 57606 3516 57612 3528
rect 55876 3512 56594 3516
rect 52457 3479 52515 3485
rect 55784 3488 56594 3512
rect 57567 3488 57612 3516
rect 55784 3484 55904 3488
rect 55784 3448 55812 3484
rect 51046 3420 55812 3448
rect 56566 3448 56594 3488
rect 57606 3476 57612 3488
rect 57664 3476 57670 3528
rect 58176 3516 58204 3556
rect 61105 3553 61117 3556
rect 61151 3553 61163 3587
rect 61105 3547 61163 3553
rect 61654 3544 61660 3596
rect 61712 3584 61718 3596
rect 97810 3584 97816 3596
rect 61712 3556 97816 3584
rect 61712 3544 61718 3556
rect 97810 3544 97816 3556
rect 97868 3544 97874 3596
rect 118068 3584 118096 3615
rect 109006 3556 118096 3584
rect 58250 3521 58256 3528
rect 57808 3488 58204 3516
rect 57808 3448 57836 3488
rect 58245 3476 58256 3521
rect 58308 3476 58314 3528
rect 58526 3476 58532 3528
rect 58584 3516 58590 3528
rect 68462 3516 68468 3528
rect 58584 3488 68468 3516
rect 58584 3476 58590 3488
rect 68462 3476 68468 3488
rect 68520 3476 68526 3528
rect 70762 3476 70768 3528
rect 70820 3516 70826 3528
rect 70949 3519 71007 3525
rect 70949 3516 70961 3519
rect 70820 3488 70961 3516
rect 70820 3476 70826 3488
rect 70949 3485 70961 3488
rect 70995 3485 71007 3519
rect 71590 3516 71596 3528
rect 71551 3488 71596 3516
rect 70949 3479 71007 3485
rect 71590 3476 71596 3488
rect 71648 3476 71654 3528
rect 72142 3476 72148 3528
rect 72200 3516 72206 3528
rect 72237 3519 72295 3525
rect 72237 3516 72249 3519
rect 72200 3488 72249 3516
rect 72200 3476 72206 3488
rect 72237 3485 72249 3488
rect 72283 3485 72295 3519
rect 72237 3479 72295 3485
rect 72605 3519 72663 3525
rect 72605 3485 72617 3519
rect 72651 3516 72663 3519
rect 73065 3519 73123 3525
rect 73065 3516 73077 3519
rect 72651 3488 73077 3516
rect 72651 3485 72663 3488
rect 72605 3479 72663 3485
rect 73065 3485 73077 3488
rect 73111 3516 73123 3519
rect 73154 3516 73160 3528
rect 73111 3488 73160 3516
rect 73111 3485 73123 3488
rect 73065 3479 73123 3485
rect 73154 3476 73160 3488
rect 73212 3476 73218 3528
rect 74166 3476 74172 3528
rect 74224 3516 74230 3528
rect 74224 3488 74269 3516
rect 74224 3476 74230 3488
rect 74902 3476 74908 3528
rect 74960 3516 74966 3528
rect 74997 3519 75055 3525
rect 74997 3516 75009 3519
rect 74960 3488 75009 3516
rect 74960 3476 74966 3488
rect 74997 3485 75009 3488
rect 75043 3485 75055 3519
rect 74997 3479 75055 3485
rect 76101 3519 76159 3525
rect 76101 3485 76113 3519
rect 76147 3516 76159 3519
rect 78030 3516 78036 3528
rect 76147 3488 78036 3516
rect 76147 3485 76159 3488
rect 76101 3479 76159 3485
rect 78030 3476 78036 3488
rect 78088 3476 78094 3528
rect 58245 3475 58303 3476
rect 59538 3448 59544 3460
rect 56566 3420 57836 3448
rect 59499 3420 59544 3448
rect 47360 3408 47366 3420
rect 59538 3408 59544 3420
rect 59596 3408 59602 3460
rect 60274 3408 60280 3460
rect 60332 3448 60338 3460
rect 60921 3451 60979 3457
rect 60921 3448 60933 3451
rect 60332 3420 60933 3448
rect 60332 3408 60338 3420
rect 60921 3417 60933 3420
rect 60967 3417 60979 3451
rect 60921 3411 60979 3417
rect 66990 3408 66996 3460
rect 67048 3448 67054 3460
rect 101490 3448 101496 3460
rect 67048 3420 101496 3448
rect 67048 3408 67054 3420
rect 101490 3408 101496 3420
rect 101548 3408 101554 3460
rect 1302 3340 1308 3392
rect 1360 3380 1366 3392
rect 2041 3383 2099 3389
rect 2041 3380 2053 3383
rect 1360 3352 2053 3380
rect 1360 3340 1366 3352
rect 2041 3349 2053 3352
rect 2087 3349 2099 3383
rect 2041 3343 2099 3349
rect 2685 3383 2743 3389
rect 2685 3349 2697 3383
rect 2731 3380 2743 3383
rect 2866 3380 2872 3392
rect 2731 3352 2872 3380
rect 2731 3349 2743 3352
rect 2685 3343 2743 3349
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 32677 3383 32735 3389
rect 32677 3349 32689 3383
rect 32723 3380 32735 3383
rect 41782 3380 41788 3392
rect 32723 3352 41788 3380
rect 32723 3349 32735 3352
rect 32677 3343 32735 3349
rect 41782 3340 41788 3352
rect 41840 3340 41846 3392
rect 42426 3340 42432 3392
rect 42484 3380 42490 3392
rect 42613 3383 42671 3389
rect 42613 3380 42625 3383
rect 42484 3352 42625 3380
rect 42484 3340 42490 3352
rect 42613 3349 42625 3352
rect 42659 3349 42671 3383
rect 42613 3343 42671 3349
rect 42794 3340 42800 3392
rect 42852 3340 42858 3392
rect 45830 3380 45836 3392
rect 45791 3352 45836 3380
rect 45830 3340 45836 3352
rect 45888 3340 45894 3392
rect 46842 3380 46848 3392
rect 46803 3352 46848 3380
rect 46842 3340 46848 3352
rect 46900 3340 46906 3392
rect 47486 3380 47492 3392
rect 47447 3352 47492 3380
rect 47486 3340 47492 3352
rect 47544 3340 47550 3392
rect 47578 3340 47584 3392
rect 47636 3380 47642 3392
rect 50798 3380 50804 3392
rect 47636 3352 50804 3380
rect 47636 3340 47642 3352
rect 50798 3340 50804 3352
rect 50856 3340 50862 3392
rect 50890 3340 50896 3392
rect 50948 3380 50954 3392
rect 57146 3380 57152 3392
rect 50948 3352 57152 3380
rect 50948 3340 50954 3352
rect 57146 3340 57152 3352
rect 57204 3340 57210 3392
rect 57330 3340 57336 3392
rect 57388 3380 57394 3392
rect 57425 3383 57483 3389
rect 57425 3380 57437 3383
rect 57388 3352 57437 3380
rect 57388 3340 57394 3352
rect 57425 3349 57437 3352
rect 57471 3349 57483 3383
rect 57425 3343 57483 3349
rect 58069 3383 58127 3389
rect 58069 3349 58081 3383
rect 58115 3380 58127 3383
rect 58158 3380 58164 3392
rect 58115 3352 58164 3380
rect 58115 3349 58127 3352
rect 58069 3343 58127 3349
rect 58158 3340 58164 3352
rect 58216 3340 58222 3392
rect 70210 3340 70216 3392
rect 70268 3380 70274 3392
rect 70765 3383 70823 3389
rect 70765 3380 70777 3383
rect 70268 3352 70777 3380
rect 70268 3340 70274 3352
rect 70765 3349 70777 3352
rect 70811 3349 70823 3383
rect 70765 3343 70823 3349
rect 70854 3340 70860 3392
rect 70912 3380 70918 3392
rect 71409 3383 71467 3389
rect 71409 3380 71421 3383
rect 70912 3352 71421 3380
rect 70912 3340 70918 3352
rect 71409 3349 71421 3352
rect 71455 3349 71467 3383
rect 72050 3380 72056 3392
rect 72011 3352 72056 3380
rect 71409 3343 71467 3349
rect 72050 3340 72056 3352
rect 72108 3340 72114 3392
rect 72881 3383 72939 3389
rect 72881 3349 72893 3383
rect 72927 3380 72939 3383
rect 74166 3380 74172 3392
rect 72927 3352 74172 3380
rect 72927 3349 72939 3352
rect 72881 3343 72939 3349
rect 74166 3340 74172 3352
rect 74224 3340 74230 3392
rect 74534 3340 74540 3392
rect 74592 3380 74598 3392
rect 74813 3383 74871 3389
rect 74813 3380 74825 3383
rect 74592 3352 74825 3380
rect 74592 3340 74598 3352
rect 74813 3349 74825 3352
rect 74859 3349 74871 3383
rect 74813 3343 74871 3349
rect 75454 3340 75460 3392
rect 75512 3380 75518 3392
rect 75917 3383 75975 3389
rect 75917 3380 75929 3383
rect 75512 3352 75929 3380
rect 75512 3340 75518 3352
rect 75917 3349 75929 3352
rect 75963 3349 75975 3383
rect 75917 3343 75975 3349
rect 76006 3340 76012 3392
rect 76064 3380 76070 3392
rect 77110 3380 77116 3392
rect 76064 3352 77116 3380
rect 76064 3340 76070 3352
rect 77110 3340 77116 3352
rect 77168 3340 77174 3392
rect 77478 3340 77484 3392
rect 77536 3380 77542 3392
rect 109006 3380 109034 3556
rect 116581 3519 116639 3525
rect 116581 3485 116593 3519
rect 116627 3516 116639 3519
rect 117406 3516 117412 3528
rect 116627 3488 117268 3516
rect 117367 3488 117412 3516
rect 116627 3485 116639 3488
rect 116581 3479 116639 3485
rect 77536 3352 109034 3380
rect 116397 3383 116455 3389
rect 77536 3340 77542 3352
rect 116397 3349 116409 3383
rect 116443 3380 116455 3383
rect 116670 3380 116676 3392
rect 116443 3352 116676 3380
rect 116443 3349 116455 3352
rect 116397 3343 116455 3349
rect 116670 3340 116676 3352
rect 116728 3340 116734 3392
rect 117240 3389 117268 3488
rect 117406 3476 117412 3488
rect 117464 3476 117470 3528
rect 117866 3516 117872 3528
rect 117827 3488 117872 3516
rect 117866 3476 117872 3488
rect 117924 3476 117930 3528
rect 117225 3383 117283 3389
rect 117225 3349 117237 3383
rect 117271 3349 117283 3383
rect 117225 3343 117283 3349
rect 1104 3290 118864 3312
rect 1104 3238 30398 3290
rect 30450 3238 30462 3290
rect 30514 3238 30526 3290
rect 30578 3238 30590 3290
rect 30642 3238 30654 3290
rect 30706 3238 59846 3290
rect 59898 3238 59910 3290
rect 59962 3238 59974 3290
rect 60026 3238 60038 3290
rect 60090 3238 60102 3290
rect 60154 3238 89294 3290
rect 89346 3238 89358 3290
rect 89410 3238 89422 3290
rect 89474 3238 89486 3290
rect 89538 3238 89550 3290
rect 89602 3238 118864 3290
rect 1104 3216 118864 3238
rect 2130 3176 2136 3188
rect 2091 3148 2136 3176
rect 2130 3136 2136 3148
rect 2188 3136 2194 3188
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 2590 3136 2596 3188
rect 2648 3176 2654 3188
rect 2648 3148 6914 3176
rect 2648 3136 2654 3148
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3108 1915 3111
rect 2774 3108 2780 3120
rect 1903 3080 2780 3108
rect 1903 3077 1915 3080
rect 1857 3071 1915 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 6886 3108 6914 3148
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10321 3179 10379 3185
rect 10321 3176 10333 3179
rect 10284 3148 10333 3176
rect 10284 3136 10290 3148
rect 10321 3145 10333 3148
rect 10367 3145 10379 3179
rect 20714 3176 20720 3188
rect 20675 3148 20720 3176
rect 10321 3139 10379 3145
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 24486 3136 24492 3188
rect 24544 3176 24550 3188
rect 28902 3176 28908 3188
rect 24544 3148 28764 3176
rect 28863 3148 28908 3176
rect 24544 3136 24550 3148
rect 6886 3080 28396 3108
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 2685 3043 2743 3049
rect 2685 3040 2697 3043
rect 2648 3012 2697 3040
rect 2648 3000 2654 3012
rect 2685 3009 2697 3012
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 3510 3040 3516 3052
rect 3099 3012 3516 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 5442 3040 5448 3052
rect 5403 3012 5448 3040
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6595 3012 6929 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 6917 3009 6929 3012
rect 6963 3040 6975 3043
rect 7190 3040 7196 3052
rect 6963 3012 7196 3040
rect 6963 3009 6975 3012
rect 6917 3003 6975 3009
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 7834 3040 7840 3052
rect 7795 3012 7840 3040
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3040 10287 3043
rect 12253 3043 12311 3049
rect 12253 3040 12265 3043
rect 10275 3012 12265 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 12253 3009 12265 3012
rect 12299 3040 12311 3043
rect 12342 3040 12348 3052
rect 12299 3012 12348 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 14240 3012 14473 3040
rect 14240 3000 14246 3012
rect 14461 3009 14473 3012
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 20901 3043 20959 3049
rect 20901 3040 20913 3043
rect 20680 3012 20913 3040
rect 20680 3000 20686 3012
rect 20901 3009 20913 3012
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 23106 3000 23112 3052
rect 23164 3040 23170 3052
rect 24486 3040 24492 3052
rect 23164 3012 24492 3040
rect 23164 3000 23170 3012
rect 24486 3000 24492 3012
rect 24544 3000 24550 3052
rect 27614 3040 27620 3052
rect 27575 3012 27620 3040
rect 27614 3000 27620 3012
rect 27672 3000 27678 3052
rect 28261 3043 28319 3049
rect 28261 3009 28273 3043
rect 28307 3009 28319 3043
rect 28261 3003 28319 3009
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 7742 2972 7748 2984
rect 7607 2944 7748 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 28276 2972 28304 3003
rect 27448 2944 28304 2972
rect 28368 2972 28396 3080
rect 28736 3049 28764 3148
rect 28902 3136 28908 3148
rect 28960 3136 28966 3188
rect 29638 3176 29644 3188
rect 29599 3148 29644 3176
rect 29638 3136 29644 3148
rect 29696 3136 29702 3188
rect 41230 3176 41236 3188
rect 31726 3148 41236 3176
rect 31726 3108 31754 3148
rect 41230 3136 41236 3148
rect 41288 3136 41294 3188
rect 41693 3179 41751 3185
rect 41693 3145 41705 3179
rect 41739 3145 41751 3179
rect 41693 3139 41751 3145
rect 32950 3108 32956 3120
rect 28828 3080 31754 3108
rect 32911 3080 32956 3108
rect 28721 3043 28779 3049
rect 28721 3009 28733 3043
rect 28767 3009 28779 3043
rect 28721 3003 28779 3009
rect 28828 2972 28856 3080
rect 32950 3068 32956 3080
rect 33008 3068 33014 3120
rect 37568 3080 38424 3108
rect 28902 3000 28908 3052
rect 28960 3040 28966 3052
rect 29549 3043 29607 3049
rect 29549 3040 29561 3043
rect 28960 3012 29561 3040
rect 28960 3000 28966 3012
rect 29549 3009 29561 3012
rect 29595 3009 29607 3043
rect 29549 3003 29607 3009
rect 31573 3043 31631 3049
rect 31573 3009 31585 3043
rect 31619 3040 31631 3043
rect 32585 3043 32643 3049
rect 32585 3040 32597 3043
rect 31619 3012 32597 3040
rect 31619 3009 31631 3012
rect 31573 3003 31631 3009
rect 28368 2944 28856 2972
rect 14 2864 20 2916
rect 72 2904 78 2916
rect 27448 2913 27476 2944
rect 3329 2907 3387 2913
rect 3329 2904 3341 2907
rect 72 2876 3341 2904
rect 72 2864 78 2876
rect 3329 2873 3341 2876
rect 3375 2873 3387 2907
rect 3329 2867 3387 2873
rect 14277 2907 14335 2913
rect 14277 2873 14289 2907
rect 14323 2904 14335 2907
rect 27433 2907 27491 2913
rect 14323 2876 27384 2904
rect 14323 2873 14335 2876
rect 14277 2867 14335 2873
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5261 2839 5319 2845
rect 5261 2836 5273 2839
rect 5224 2808 5273 2836
rect 5224 2796 5230 2808
rect 5261 2805 5273 2808
rect 5307 2805 5319 2839
rect 5261 2799 5319 2805
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 5868 2808 6377 2836
rect 5868 2796 5874 2808
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 6365 2799 6423 2805
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 7193 2839 7251 2845
rect 7193 2836 7205 2839
rect 7156 2808 7205 2836
rect 7156 2796 7162 2808
rect 7193 2805 7205 2808
rect 7239 2805 7251 2839
rect 7193 2799 7251 2805
rect 12069 2839 12127 2845
rect 12069 2805 12081 2839
rect 12115 2836 12127 2839
rect 12618 2836 12624 2848
rect 12115 2808 12624 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 24305 2839 24363 2845
rect 24305 2805 24317 2839
rect 24351 2836 24363 2839
rect 24762 2836 24768 2848
rect 24351 2808 24768 2836
rect 24351 2805 24363 2808
rect 24305 2799 24363 2805
rect 24762 2796 24768 2808
rect 24820 2796 24826 2848
rect 26418 2836 26424 2848
rect 26379 2808 26424 2836
rect 26418 2796 26424 2808
rect 26476 2796 26482 2848
rect 27356 2836 27384 2876
rect 27433 2873 27445 2907
rect 27479 2873 27491 2907
rect 31726 2904 31754 3012
rect 32585 3009 32597 3012
rect 32631 3009 32643 3043
rect 33594 3040 33600 3052
rect 33555 3012 33600 3040
rect 32585 3003 32643 3009
rect 33594 3000 33600 3012
rect 33652 3000 33658 3052
rect 34790 3000 34796 3052
rect 34848 3040 34854 3052
rect 35069 3043 35127 3049
rect 35069 3040 35081 3043
rect 34848 3012 35081 3040
rect 34848 3000 34854 3012
rect 35069 3009 35081 3012
rect 35115 3009 35127 3043
rect 35069 3003 35127 3009
rect 35434 3000 35440 3052
rect 35492 3040 35498 3052
rect 35529 3043 35587 3049
rect 35529 3040 35541 3043
rect 35492 3012 35541 3040
rect 35492 3000 35498 3012
rect 35529 3009 35541 3012
rect 35575 3009 35587 3043
rect 35529 3003 35587 3009
rect 36078 3000 36084 3052
rect 36136 3040 36142 3052
rect 36449 3043 36507 3049
rect 36449 3040 36461 3043
rect 36136 3012 36461 3040
rect 36136 3000 36142 3012
rect 36449 3009 36461 3012
rect 36495 3009 36507 3043
rect 36449 3003 36507 3009
rect 37568 2972 37596 3080
rect 37642 3000 37648 3052
rect 37700 3040 37706 3052
rect 38289 3043 38347 3049
rect 37700 3012 37745 3040
rect 37700 3000 37706 3012
rect 38289 3009 38301 3043
rect 38335 3009 38347 3043
rect 38289 3003 38347 3009
rect 37734 2972 37740 2984
rect 34900 2944 37596 2972
rect 37695 2944 37740 2972
rect 34900 2913 34928 2944
rect 37734 2932 37740 2944
rect 37792 2932 37798 2984
rect 37826 2932 37832 2984
rect 37884 2972 37890 2984
rect 37884 2944 37929 2972
rect 37884 2932 37890 2944
rect 27433 2867 27491 2873
rect 28000 2876 31754 2904
rect 34885 2907 34943 2913
rect 28000 2836 28028 2876
rect 34885 2873 34897 2907
rect 34931 2873 34943 2907
rect 35710 2904 35716 2916
rect 35671 2876 35716 2904
rect 34885 2867 34943 2873
rect 35710 2864 35716 2876
rect 35768 2864 35774 2916
rect 37277 2907 37335 2913
rect 37277 2873 37289 2907
rect 37323 2904 37335 2907
rect 38304 2904 38332 3003
rect 37323 2876 38332 2904
rect 38396 2904 38424 3080
rect 41708 3052 41736 3139
rect 41782 3136 41788 3188
rect 41840 3176 41846 3188
rect 42794 3176 42800 3188
rect 41840 3148 42800 3176
rect 41840 3136 41846 3148
rect 42794 3136 42800 3148
rect 42852 3136 42858 3188
rect 43073 3179 43131 3185
rect 43073 3145 43085 3179
rect 43119 3176 43131 3179
rect 43901 3179 43959 3185
rect 43901 3176 43913 3179
rect 43119 3148 43913 3176
rect 43119 3145 43131 3148
rect 43073 3139 43131 3145
rect 43901 3145 43913 3148
rect 43947 3145 43959 3179
rect 47670 3176 47676 3188
rect 43901 3139 43959 3145
rect 45572 3148 47676 3176
rect 42978 3068 42984 3120
rect 43036 3108 43042 3120
rect 45572 3117 45600 3148
rect 47670 3136 47676 3148
rect 47728 3136 47734 3188
rect 47765 3179 47823 3185
rect 47765 3145 47777 3179
rect 47811 3145 47823 3179
rect 47765 3139 47823 3145
rect 45557 3111 45615 3117
rect 43036 3080 43081 3108
rect 43036 3068 43042 3080
rect 45557 3077 45569 3111
rect 45603 3077 45615 3111
rect 47029 3111 47087 3117
rect 45557 3071 45615 3077
rect 46032 3080 46980 3108
rect 39574 3040 39580 3052
rect 39535 3012 39580 3040
rect 39574 3000 39580 3012
rect 39632 3000 39638 3052
rect 40402 3040 40408 3052
rect 40363 3012 40408 3040
rect 40402 3000 40408 3012
rect 40460 3000 40466 3052
rect 41690 3000 41696 3052
rect 41748 3000 41754 3052
rect 41877 3043 41935 3049
rect 41877 3009 41889 3043
rect 41923 3040 41935 3043
rect 41966 3040 41972 3052
rect 41923 3012 41972 3040
rect 41923 3009 41935 3012
rect 41877 3003 41935 3009
rect 41966 3000 41972 3012
rect 42024 3000 42030 3052
rect 43806 3000 43812 3052
rect 43864 3040 43870 3052
rect 44085 3043 44143 3049
rect 44085 3040 44097 3043
rect 43864 3012 44097 3040
rect 43864 3000 43870 3012
rect 44085 3009 44097 3012
rect 44131 3009 44143 3043
rect 44085 3003 44143 3009
rect 45370 3000 45376 3052
rect 45428 3040 45434 3052
rect 46032 3049 46060 3080
rect 46017 3043 46075 3049
rect 45428 3012 45473 3040
rect 45428 3000 45434 3012
rect 46017 3009 46029 3043
rect 46063 3009 46075 3043
rect 46017 3003 46075 3009
rect 46382 3000 46388 3052
rect 46440 3040 46446 3052
rect 46845 3043 46903 3049
rect 46845 3040 46857 3043
rect 46440 3012 46857 3040
rect 46440 3000 46446 3012
rect 46845 3009 46857 3012
rect 46891 3009 46903 3043
rect 46952 3040 46980 3080
rect 47029 3077 47041 3111
rect 47075 3108 47087 3111
rect 47118 3108 47124 3120
rect 47075 3080 47124 3108
rect 47075 3077 47087 3080
rect 47029 3071 47087 3077
rect 47118 3068 47124 3080
rect 47176 3068 47182 3120
rect 47780 3108 47808 3139
rect 47854 3136 47860 3188
rect 47912 3176 47918 3188
rect 57606 3176 57612 3188
rect 47912 3148 57612 3176
rect 47912 3136 47918 3148
rect 57606 3136 57612 3148
rect 57664 3136 57670 3188
rect 58066 3176 58072 3188
rect 58027 3148 58072 3176
rect 58066 3136 58072 3148
rect 58124 3136 58130 3188
rect 76006 3176 76012 3188
rect 58176 3148 76012 3176
rect 47780 3080 48636 3108
rect 47578 3040 47584 3052
rect 46952 3012 47584 3040
rect 46845 3003 46903 3009
rect 47578 3000 47584 3012
rect 47636 3000 47642 3052
rect 47946 3040 47952 3052
rect 47907 3012 47952 3040
rect 47946 3000 47952 3012
rect 48004 3000 48010 3052
rect 48608 3049 48636 3080
rect 48700 3080 54064 3108
rect 48593 3043 48651 3049
rect 48593 3009 48605 3043
rect 48639 3009 48651 3043
rect 48593 3003 48651 3009
rect 40218 2932 40224 2984
rect 40276 2972 40282 2984
rect 40497 2975 40555 2981
rect 40497 2972 40509 2975
rect 40276 2944 40509 2972
rect 40276 2932 40282 2944
rect 40497 2941 40509 2944
rect 40543 2941 40555 2975
rect 40678 2972 40684 2984
rect 40639 2944 40684 2972
rect 40497 2935 40555 2941
rect 40678 2932 40684 2944
rect 40736 2932 40742 2984
rect 43254 2972 43260 2984
rect 41616 2944 43116 2972
rect 43215 2944 43260 2972
rect 41616 2904 41644 2944
rect 38396 2876 41644 2904
rect 43088 2904 43116 2944
rect 43254 2932 43260 2944
rect 43312 2932 43318 2984
rect 45830 2932 45836 2984
rect 45888 2972 45894 2984
rect 48700 2972 48728 3080
rect 51166 3040 51172 3052
rect 51127 3012 51172 3040
rect 51166 3000 51172 3012
rect 51224 3000 51230 3052
rect 51905 3043 51963 3049
rect 51905 3009 51917 3043
rect 51951 3040 51963 3043
rect 52730 3040 52736 3052
rect 51951 3012 52736 3040
rect 51951 3009 51963 3012
rect 51905 3003 51963 3009
rect 52730 3000 52736 3012
rect 52788 3000 52794 3052
rect 52822 3000 52828 3052
rect 52880 3040 52886 3052
rect 53101 3043 53159 3049
rect 53101 3040 53113 3043
rect 52880 3012 53113 3040
rect 52880 3000 52886 3012
rect 53101 3009 53113 3012
rect 53147 3009 53159 3043
rect 54036 3040 54064 3080
rect 54110 3068 54116 3120
rect 54168 3108 54174 3120
rect 56686 3108 56692 3120
rect 54168 3080 56692 3108
rect 54168 3068 54174 3080
rect 56686 3068 56692 3080
rect 56744 3068 56750 3120
rect 56962 3108 56968 3120
rect 56923 3080 56968 3108
rect 56962 3068 56968 3080
rect 57020 3068 57026 3120
rect 57057 3111 57115 3117
rect 57057 3077 57069 3111
rect 57103 3108 57115 3111
rect 57146 3108 57152 3120
rect 57103 3080 57152 3108
rect 57103 3077 57115 3080
rect 57057 3071 57115 3077
rect 57146 3068 57152 3080
rect 57204 3068 57210 3120
rect 57974 3068 57980 3120
rect 58032 3108 58038 3120
rect 58176 3108 58204 3148
rect 76006 3136 76012 3148
rect 76064 3136 76070 3188
rect 76929 3179 76987 3185
rect 76929 3176 76941 3179
rect 76760 3148 76941 3176
rect 58032 3080 58204 3108
rect 58032 3068 58038 3080
rect 59538 3068 59544 3120
rect 59596 3108 59602 3120
rect 60829 3111 60887 3117
rect 60829 3108 60841 3111
rect 59596 3080 60841 3108
rect 59596 3068 59602 3080
rect 60829 3077 60841 3080
rect 60875 3077 60887 3111
rect 60829 3071 60887 3077
rect 61013 3111 61071 3117
rect 61013 3077 61025 3111
rect 61059 3108 61071 3111
rect 61654 3108 61660 3120
rect 61059 3080 61660 3108
rect 61059 3077 61071 3080
rect 61013 3071 61071 3077
rect 61654 3068 61660 3080
rect 61712 3068 61718 3120
rect 61746 3068 61752 3120
rect 61804 3108 61810 3120
rect 70302 3108 70308 3120
rect 61804 3080 70308 3108
rect 61804 3068 61810 3080
rect 70302 3068 70308 3080
rect 70360 3068 70366 3120
rect 70578 3108 70584 3120
rect 70539 3080 70584 3108
rect 70578 3068 70584 3080
rect 70636 3068 70642 3120
rect 74534 3108 74540 3120
rect 74495 3080 74540 3108
rect 74534 3068 74540 3080
rect 74592 3108 74598 3120
rect 75273 3111 75331 3117
rect 75273 3108 75285 3111
rect 74592 3080 75285 3108
rect 74592 3068 74598 3080
rect 75273 3077 75285 3080
rect 75319 3077 75331 3111
rect 75273 3071 75331 3077
rect 75362 3068 75368 3120
rect 75420 3108 75426 3120
rect 76760 3108 76788 3148
rect 76929 3145 76941 3148
rect 76975 3145 76987 3179
rect 76929 3139 76987 3145
rect 77110 3136 77116 3188
rect 77168 3176 77174 3188
rect 85298 3176 85304 3188
rect 77168 3148 85304 3176
rect 77168 3136 77174 3148
rect 85298 3136 85304 3148
rect 85356 3136 85362 3188
rect 102778 3176 102784 3188
rect 96586 3148 102784 3176
rect 75420 3080 76788 3108
rect 75420 3068 75426 3080
rect 77018 3068 77024 3120
rect 77076 3108 77082 3120
rect 96586 3108 96614 3148
rect 102778 3136 102784 3148
rect 102836 3136 102842 3188
rect 104250 3136 104256 3188
rect 104308 3176 104314 3188
rect 117130 3176 117136 3188
rect 104308 3148 116992 3176
rect 117091 3148 117136 3176
rect 104308 3136 104314 3148
rect 77076 3080 96614 3108
rect 101309 3111 101367 3117
rect 77076 3068 77082 3080
rect 101309 3077 101321 3111
rect 101355 3108 101367 3111
rect 103974 3108 103980 3120
rect 101355 3080 103980 3108
rect 101355 3077 101367 3080
rect 101309 3071 101367 3077
rect 103974 3068 103980 3080
rect 104032 3068 104038 3120
rect 107470 3108 107476 3120
rect 107431 3080 107476 3108
rect 107470 3068 107476 3080
rect 107528 3068 107534 3120
rect 109770 3068 109776 3120
rect 109828 3108 109834 3120
rect 109828 3080 110368 3108
rect 109828 3068 109834 3080
rect 55582 3040 55588 3052
rect 54036 3012 55588 3040
rect 53101 3003 53159 3009
rect 55582 3000 55588 3012
rect 55640 3000 55646 3052
rect 55677 3043 55735 3049
rect 55677 3009 55689 3043
rect 55723 3040 55735 3043
rect 57698 3040 57704 3052
rect 55723 3012 57704 3040
rect 55723 3009 55735 3012
rect 55677 3003 55735 3009
rect 57698 3000 57704 3012
rect 57756 3000 57762 3052
rect 57873 3043 57931 3049
rect 57873 3040 57885 3043
rect 57808 3012 57885 3040
rect 45888 2944 48728 2972
rect 45888 2932 45894 2944
rect 50614 2932 50620 2984
rect 50672 2972 50678 2984
rect 57241 2975 57299 2981
rect 50672 2944 55628 2972
rect 50672 2932 50678 2944
rect 48038 2904 48044 2916
rect 43088 2876 48044 2904
rect 37323 2873 37335 2876
rect 37277 2867 37335 2873
rect 48038 2864 48044 2876
rect 48096 2864 48102 2916
rect 52089 2907 52147 2913
rect 52089 2904 52101 2907
rect 48148 2876 52101 2904
rect 27356 2808 28028 2836
rect 28077 2839 28135 2845
rect 28077 2805 28089 2839
rect 28123 2836 28135 2839
rect 28350 2836 28356 2848
rect 28123 2808 28356 2836
rect 28123 2805 28135 2808
rect 28077 2799 28135 2805
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 31389 2839 31447 2845
rect 31389 2805 31401 2839
rect 31435 2836 31447 2839
rect 31570 2836 31576 2848
rect 31435 2808 31576 2836
rect 31435 2805 31447 2808
rect 31389 2799 31447 2805
rect 31570 2796 31576 2808
rect 31628 2796 31634 2848
rect 32858 2796 32864 2848
rect 32916 2836 32922 2848
rect 33413 2839 33471 2845
rect 33413 2836 33425 2839
rect 32916 2808 33425 2836
rect 32916 2796 32922 2808
rect 33413 2805 33425 2808
rect 33459 2805 33471 2839
rect 36262 2836 36268 2848
rect 36223 2808 36268 2836
rect 33413 2799 33471 2805
rect 36262 2796 36268 2808
rect 36320 2796 36326 2848
rect 37642 2796 37648 2848
rect 37700 2836 37706 2848
rect 38105 2839 38163 2845
rect 38105 2836 38117 2839
rect 37700 2808 38117 2836
rect 37700 2796 37706 2808
rect 38105 2805 38117 2808
rect 38151 2805 38163 2839
rect 39390 2836 39396 2848
rect 39351 2808 39396 2836
rect 38105 2799 38163 2805
rect 39390 2796 39396 2808
rect 39448 2796 39454 2848
rect 40034 2836 40040 2848
rect 39995 2808 40040 2836
rect 40034 2796 40040 2808
rect 40092 2796 40098 2848
rect 42610 2836 42616 2848
rect 42571 2808 42616 2836
rect 42610 2796 42616 2808
rect 42668 2796 42674 2848
rect 46198 2836 46204 2848
rect 46159 2808 46204 2836
rect 46198 2796 46204 2808
rect 46256 2796 46262 2848
rect 46290 2796 46296 2848
rect 46348 2836 46354 2848
rect 48148 2836 48176 2876
rect 52089 2873 52101 2876
rect 52135 2873 52147 2907
rect 55600 2904 55628 2944
rect 57241 2941 57253 2975
rect 57287 2972 57299 2975
rect 57422 2972 57428 2984
rect 57287 2944 57428 2972
rect 57287 2941 57299 2944
rect 57241 2935 57299 2941
rect 57422 2932 57428 2944
rect 57480 2932 57486 2984
rect 57808 2972 57836 3012
rect 57873 3009 57885 3012
rect 57919 3009 57931 3043
rect 57873 3003 57931 3009
rect 58989 3043 59047 3049
rect 58989 3009 59001 3043
rect 59035 3040 59047 3043
rect 59722 3040 59728 3052
rect 59035 3012 59584 3040
rect 59683 3012 59728 3040
rect 59035 3009 59047 3012
rect 58989 3003 59047 3009
rect 57974 2972 57980 2984
rect 57808 2944 57980 2972
rect 57974 2932 57980 2944
rect 58032 2932 58038 2984
rect 59446 2972 59452 2984
rect 59407 2944 59452 2972
rect 59446 2932 59452 2944
rect 59504 2932 59510 2984
rect 59556 2972 59584 3012
rect 59722 3000 59728 3012
rect 59780 3000 59786 3052
rect 61838 3000 61844 3052
rect 61896 3040 61902 3052
rect 62117 3043 62175 3049
rect 62117 3040 62129 3043
rect 61896 3012 62129 3040
rect 61896 3000 61902 3012
rect 62117 3009 62129 3012
rect 62163 3009 62175 3043
rect 62117 3003 62175 3009
rect 64046 3000 64052 3052
rect 64104 3040 64110 3052
rect 64417 3043 64475 3049
rect 64417 3040 64429 3043
rect 64104 3012 64429 3040
rect 64104 3000 64110 3012
rect 64417 3009 64429 3012
rect 64463 3009 64475 3043
rect 64417 3003 64475 3009
rect 64506 3000 64512 3052
rect 64564 3040 64570 3052
rect 65245 3043 65303 3049
rect 65245 3040 65257 3043
rect 64564 3012 65257 3040
rect 64564 3000 64570 3012
rect 65245 3009 65257 3012
rect 65291 3009 65303 3043
rect 65245 3003 65303 3009
rect 66349 3043 66407 3049
rect 66349 3009 66361 3043
rect 66395 3040 66407 3043
rect 66714 3040 66720 3052
rect 66395 3012 66720 3040
rect 66395 3009 66407 3012
rect 66349 3003 66407 3009
rect 66714 3000 66720 3012
rect 66772 3000 66778 3052
rect 66990 3040 66996 3052
rect 66951 3012 66996 3040
rect 66990 3000 66996 3012
rect 67048 3000 67054 3052
rect 68278 3000 68284 3052
rect 68336 3040 68342 3052
rect 68557 3043 68615 3049
rect 68557 3040 68569 3043
rect 68336 3012 68569 3040
rect 68336 3000 68342 3012
rect 68557 3009 68569 3012
rect 68603 3009 68615 3043
rect 68557 3003 68615 3009
rect 69566 3000 69572 3052
rect 69624 3040 69630 3052
rect 69845 3043 69903 3049
rect 69845 3040 69857 3043
rect 69624 3012 69857 3040
rect 69624 3000 69630 3012
rect 69845 3009 69857 3012
rect 69891 3009 69903 3043
rect 69845 3003 69903 3009
rect 70394 3000 70400 3052
rect 70452 3040 70458 3052
rect 71225 3044 71283 3049
rect 71314 3044 71320 3052
rect 71225 3043 71320 3044
rect 70452 3012 70497 3040
rect 70780 3012 70992 3040
rect 70452 3000 70458 3012
rect 59998 2972 60004 2984
rect 59556 2944 60004 2972
rect 59998 2932 60004 2944
rect 60056 2932 60062 2984
rect 69934 2932 69940 2984
rect 69992 2972 69998 2984
rect 70780 2972 70808 3012
rect 69992 2944 70808 2972
rect 70964 2972 70992 3012
rect 71225 3009 71237 3043
rect 71271 3016 71320 3043
rect 71271 3009 71283 3016
rect 71225 3003 71283 3009
rect 71314 3000 71320 3016
rect 71372 3000 71378 3052
rect 72234 3040 72240 3052
rect 72195 3012 72240 3040
rect 72234 3000 72240 3012
rect 72292 3000 72298 3052
rect 72326 3000 72332 3052
rect 72384 3040 72390 3052
rect 73525 3043 73583 3049
rect 73525 3040 73537 3043
rect 72384 3012 72429 3040
rect 72528 3012 73537 3040
rect 72384 3000 72390 3012
rect 72421 2975 72479 2981
rect 72421 2972 72433 2975
rect 70964 2944 72433 2972
rect 69992 2932 69998 2944
rect 72421 2941 72433 2944
rect 72467 2941 72479 2975
rect 72421 2935 72479 2941
rect 64598 2904 64604 2916
rect 55600 2876 58940 2904
rect 64559 2876 64604 2904
rect 52089 2867 52147 2873
rect 46348 2808 48176 2836
rect 46348 2796 46354 2808
rect 48314 2796 48320 2848
rect 48372 2836 48378 2848
rect 48409 2839 48467 2845
rect 48409 2836 48421 2839
rect 48372 2808 48421 2836
rect 48372 2796 48378 2808
rect 48409 2805 48421 2808
rect 48455 2805 48467 2839
rect 48409 2799 48467 2805
rect 50890 2796 50896 2848
rect 50948 2836 50954 2848
rect 50985 2839 51043 2845
rect 50985 2836 50997 2839
rect 50948 2808 50997 2836
rect 50948 2796 50954 2808
rect 50985 2805 50997 2808
rect 51031 2805 51043 2839
rect 52914 2836 52920 2848
rect 52875 2808 52920 2836
rect 50985 2799 51043 2805
rect 52914 2796 52920 2808
rect 52972 2796 52978 2848
rect 55398 2796 55404 2848
rect 55456 2836 55462 2848
rect 55493 2839 55551 2845
rect 55493 2836 55505 2839
rect 55456 2808 55505 2836
rect 55456 2796 55462 2808
rect 55493 2805 55505 2808
rect 55539 2805 55551 2839
rect 55493 2799 55551 2805
rect 55858 2796 55864 2848
rect 55916 2836 55922 2848
rect 56597 2839 56655 2845
rect 56597 2836 56609 2839
rect 55916 2808 56609 2836
rect 55916 2796 55922 2808
rect 56597 2805 56609 2808
rect 56643 2805 56655 2839
rect 56597 2799 56655 2805
rect 56686 2796 56692 2848
rect 56744 2836 56750 2848
rect 57974 2836 57980 2848
rect 56744 2808 57980 2836
rect 56744 2796 56750 2808
rect 57974 2796 57980 2808
rect 58032 2796 58038 2848
rect 58066 2796 58072 2848
rect 58124 2836 58130 2848
rect 58250 2836 58256 2848
rect 58124 2808 58256 2836
rect 58124 2796 58130 2808
rect 58250 2796 58256 2808
rect 58308 2796 58314 2848
rect 58802 2836 58808 2848
rect 58763 2808 58808 2836
rect 58802 2796 58808 2808
rect 58860 2796 58866 2848
rect 58912 2836 58940 2876
rect 64598 2864 64604 2876
rect 64656 2864 64662 2916
rect 66162 2904 66168 2916
rect 66123 2876 66168 2904
rect 66162 2864 66168 2876
rect 66220 2864 66226 2916
rect 68462 2864 68468 2916
rect 68520 2904 68526 2916
rect 68520 2876 71176 2904
rect 68520 2864 68526 2876
rect 61746 2836 61752 2848
rect 58912 2808 61752 2836
rect 61746 2796 61752 2808
rect 61804 2796 61810 2848
rect 61930 2836 61936 2848
rect 61891 2808 61936 2836
rect 61930 2796 61936 2808
rect 61988 2796 61994 2848
rect 63494 2796 63500 2848
rect 63552 2836 63558 2848
rect 65061 2839 65119 2845
rect 65061 2836 65073 2839
rect 63552 2808 65073 2836
rect 63552 2796 63558 2808
rect 65061 2805 65073 2808
rect 65107 2805 65119 2839
rect 65061 2799 65119 2805
rect 66346 2796 66352 2848
rect 66404 2836 66410 2848
rect 66809 2839 66867 2845
rect 66809 2836 66821 2839
rect 66404 2808 66821 2836
rect 66404 2796 66410 2808
rect 66809 2805 66821 2808
rect 66855 2805 66867 2839
rect 66809 2799 66867 2805
rect 68094 2796 68100 2848
rect 68152 2836 68158 2848
rect 68373 2839 68431 2845
rect 68373 2836 68385 2839
rect 68152 2808 68385 2836
rect 68152 2796 68158 2808
rect 68373 2805 68385 2808
rect 68419 2805 68431 2839
rect 69658 2836 69664 2848
rect 69619 2808 69664 2836
rect 68373 2799 68431 2805
rect 69658 2796 69664 2808
rect 69716 2796 69722 2848
rect 71148 2836 71176 2876
rect 71222 2864 71228 2916
rect 71280 2904 71286 2916
rect 72326 2904 72332 2916
rect 71280 2876 72332 2904
rect 71280 2864 71286 2876
rect 72326 2864 72332 2876
rect 72384 2864 72390 2916
rect 71317 2839 71375 2845
rect 71317 2836 71329 2839
rect 71148 2808 71329 2836
rect 71317 2805 71329 2808
rect 71363 2805 71375 2839
rect 71317 2799 71375 2805
rect 71869 2839 71927 2845
rect 71869 2805 71881 2839
rect 71915 2836 71927 2839
rect 72528 2836 72556 3012
rect 73525 3009 73537 3012
rect 73571 3009 73583 3043
rect 73525 3003 73583 3009
rect 76834 3000 76840 3052
rect 76892 3040 76898 3052
rect 76892 3012 76937 3040
rect 76892 3000 76898 3012
rect 77294 3000 77300 3052
rect 77352 3040 77358 3052
rect 77849 3043 77907 3049
rect 77849 3040 77861 3043
rect 77352 3012 77861 3040
rect 77352 3000 77358 3012
rect 77849 3009 77861 3012
rect 77895 3009 77907 3043
rect 77849 3003 77907 3009
rect 80698 3000 80704 3052
rect 80756 3040 80762 3052
rect 81437 3043 81495 3049
rect 81437 3040 81449 3043
rect 80756 3012 81449 3040
rect 80756 3000 80762 3012
rect 81437 3009 81449 3012
rect 81483 3009 81495 3043
rect 87230 3040 87236 3052
rect 87191 3012 87236 3040
rect 81437 3003 81495 3009
rect 87230 3000 87236 3012
rect 87288 3000 87294 3052
rect 101490 3040 101496 3052
rect 101451 3012 101496 3040
rect 101490 3000 101496 3012
rect 101548 3000 101554 3052
rect 102686 3040 102692 3052
rect 102647 3012 102692 3040
rect 102686 3000 102692 3012
rect 102744 3000 102750 3052
rect 102778 3000 102784 3052
rect 102836 3040 102842 3052
rect 110230 3040 110236 3052
rect 102836 3012 110236 3040
rect 102836 3000 102842 3012
rect 110230 3000 110236 3012
rect 110288 3000 110294 3052
rect 110340 3049 110368 3080
rect 110325 3043 110383 3049
rect 110325 3009 110337 3043
rect 110371 3009 110383 3043
rect 110325 3003 110383 3009
rect 111426 3000 111432 3052
rect 111484 3040 111490 3052
rect 111521 3043 111579 3049
rect 111521 3040 111533 3043
rect 111484 3012 111533 3040
rect 111484 3000 111490 3012
rect 111521 3009 111533 3012
rect 111567 3009 111579 3043
rect 116210 3040 116216 3052
rect 116171 3012 116216 3040
rect 111521 3003 111579 3009
rect 116210 3000 116216 3012
rect 116268 3000 116274 3052
rect 116964 3040 116992 3148
rect 117130 3136 117136 3148
rect 117188 3136 117194 3188
rect 117041 3111 117099 3117
rect 117041 3077 117053 3111
rect 117087 3108 117099 3111
rect 118510 3108 118516 3120
rect 117087 3080 118516 3108
rect 117087 3077 117099 3080
rect 117041 3071 117099 3077
rect 118510 3068 118516 3080
rect 118568 3068 118574 3120
rect 117406 3040 117412 3052
rect 116964 3012 117412 3040
rect 117406 3000 117412 3012
rect 117464 3000 117470 3052
rect 117774 3040 117780 3052
rect 117735 3012 117780 3040
rect 117774 3000 117780 3012
rect 117832 3000 117838 3052
rect 73356 2944 76788 2972
rect 73356 2913 73384 2944
rect 73341 2907 73399 2913
rect 73341 2873 73353 2907
rect 73387 2873 73399 2907
rect 73341 2867 73399 2873
rect 75086 2864 75092 2916
rect 75144 2904 75150 2916
rect 75730 2904 75736 2916
rect 75144 2876 75736 2904
rect 75144 2864 75150 2876
rect 75730 2864 75736 2876
rect 75788 2864 75794 2916
rect 76466 2904 76472 2916
rect 76427 2876 76472 2904
rect 76466 2864 76472 2876
rect 76524 2864 76530 2916
rect 71915 2808 72556 2836
rect 71915 2805 71927 2808
rect 71869 2799 71927 2805
rect 73430 2796 73436 2848
rect 73488 2836 73494 2848
rect 74629 2839 74687 2845
rect 74629 2836 74641 2839
rect 73488 2808 74641 2836
rect 73488 2796 73494 2808
rect 74629 2805 74641 2808
rect 74675 2805 74687 2839
rect 74629 2799 74687 2805
rect 75365 2839 75423 2845
rect 75365 2805 75377 2839
rect 75411 2836 75423 2839
rect 75546 2836 75552 2848
rect 75411 2808 75552 2836
rect 75411 2805 75423 2808
rect 75365 2799 75423 2805
rect 75546 2796 75552 2808
rect 75604 2796 75610 2848
rect 76760 2836 76788 2944
rect 76926 2932 76932 2984
rect 76984 2972 76990 2984
rect 77021 2975 77079 2981
rect 77021 2972 77033 2975
rect 76984 2944 77033 2972
rect 76984 2932 76990 2944
rect 77021 2941 77033 2944
rect 77067 2941 77079 2975
rect 77021 2935 77079 2941
rect 77110 2932 77116 2984
rect 77168 2972 77174 2984
rect 118053 2975 118111 2981
rect 118053 2972 118065 2975
rect 77168 2944 118065 2972
rect 77168 2932 77174 2944
rect 118053 2941 118065 2944
rect 118099 2941 118111 2975
rect 118053 2935 118111 2941
rect 76834 2864 76840 2916
rect 76892 2904 76898 2916
rect 77665 2907 77723 2913
rect 77665 2904 77677 2907
rect 76892 2876 77677 2904
rect 76892 2864 76898 2876
rect 77665 2873 77677 2876
rect 77711 2873 77723 2907
rect 89162 2904 89168 2916
rect 77665 2867 77723 2873
rect 80026 2876 89168 2904
rect 80026 2836 80054 2876
rect 89162 2864 89168 2876
rect 89220 2864 89226 2916
rect 107654 2904 107660 2916
rect 107615 2876 107660 2904
rect 107654 2864 107660 2876
rect 107712 2864 107718 2916
rect 109494 2864 109500 2916
rect 109552 2904 109558 2916
rect 110141 2907 110199 2913
rect 110141 2904 110153 2907
rect 109552 2876 110153 2904
rect 109552 2864 109558 2876
rect 110141 2873 110153 2876
rect 110187 2873 110199 2907
rect 110141 2867 110199 2873
rect 110230 2864 110236 2916
rect 110288 2904 110294 2916
rect 111705 2907 111763 2913
rect 111705 2904 111717 2907
rect 110288 2876 111717 2904
rect 110288 2864 110294 2876
rect 111705 2873 111717 2876
rect 111751 2873 111763 2907
rect 111705 2867 111763 2873
rect 76760 2808 80054 2836
rect 81158 2796 81164 2848
rect 81216 2836 81222 2848
rect 81253 2839 81311 2845
rect 81253 2836 81265 2839
rect 81216 2808 81265 2836
rect 81216 2796 81222 2808
rect 81253 2805 81265 2808
rect 81299 2805 81311 2839
rect 81253 2799 81311 2805
rect 86954 2796 86960 2848
rect 87012 2836 87018 2848
rect 87049 2839 87107 2845
rect 87049 2836 87061 2839
rect 87012 2808 87061 2836
rect 87012 2796 87018 2808
rect 87049 2805 87061 2808
rect 87095 2805 87107 2839
rect 87049 2799 87107 2805
rect 98546 2796 98552 2848
rect 98604 2836 98610 2848
rect 99285 2839 99343 2845
rect 99285 2836 99297 2839
rect 98604 2808 99297 2836
rect 98604 2796 98610 2808
rect 99285 2805 99297 2808
rect 99331 2805 99343 2839
rect 99285 2799 99343 2805
rect 102410 2796 102416 2848
rect 102468 2836 102474 2848
rect 102505 2839 102563 2845
rect 102505 2836 102517 2839
rect 102468 2808 102517 2836
rect 102468 2796 102474 2808
rect 102505 2805 102517 2808
rect 102551 2805 102563 2839
rect 109770 2836 109776 2848
rect 109731 2808 109776 2836
rect 102505 2799 102563 2805
rect 109770 2796 109776 2808
rect 109828 2796 109834 2848
rect 115934 2796 115940 2848
rect 115992 2836 115998 2848
rect 116029 2839 116087 2845
rect 116029 2836 116041 2839
rect 115992 2808 116041 2836
rect 115992 2796 115998 2808
rect 116029 2805 116041 2808
rect 116075 2805 116087 2839
rect 116029 2799 116087 2805
rect 1104 2746 118864 2768
rect 1104 2694 15674 2746
rect 15726 2694 15738 2746
rect 15790 2694 15802 2746
rect 15854 2694 15866 2746
rect 15918 2694 15930 2746
rect 15982 2694 45122 2746
rect 45174 2694 45186 2746
rect 45238 2694 45250 2746
rect 45302 2694 45314 2746
rect 45366 2694 45378 2746
rect 45430 2694 74570 2746
rect 74622 2694 74634 2746
rect 74686 2694 74698 2746
rect 74750 2694 74762 2746
rect 74814 2694 74826 2746
rect 74878 2694 104018 2746
rect 104070 2694 104082 2746
rect 104134 2694 104146 2746
rect 104198 2694 104210 2746
rect 104262 2694 104274 2746
rect 104326 2694 118864 2746
rect 1104 2672 118864 2694
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 14642 2632 14648 2644
rect 14603 2604 14648 2632
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 19426 2592 19432 2644
rect 19484 2632 19490 2644
rect 19797 2635 19855 2641
rect 19797 2632 19809 2635
rect 19484 2604 19809 2632
rect 19484 2592 19490 2604
rect 19797 2601 19809 2604
rect 19843 2632 19855 2635
rect 22462 2632 22468 2644
rect 19843 2604 22468 2632
rect 19843 2601 19855 2604
rect 19797 2595 19855 2601
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 22649 2635 22707 2641
rect 22649 2601 22661 2635
rect 22695 2632 22707 2635
rect 23106 2632 23112 2644
rect 22695 2604 23112 2632
rect 22695 2601 22707 2604
rect 22649 2595 22707 2601
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 23290 2632 23296 2644
rect 23251 2604 23296 2632
rect 23290 2592 23296 2604
rect 23348 2592 23354 2644
rect 25406 2632 25412 2644
rect 25367 2604 25412 2632
rect 25406 2592 25412 2604
rect 25464 2592 25470 2644
rect 26973 2635 27031 2641
rect 26973 2601 26985 2635
rect 27019 2632 27031 2635
rect 27614 2632 27620 2644
rect 27019 2604 27620 2632
rect 27019 2601 27031 2604
rect 26973 2595 27031 2601
rect 27614 2592 27620 2604
rect 27672 2592 27678 2644
rect 28810 2632 28816 2644
rect 28771 2604 28816 2632
rect 28810 2592 28816 2604
rect 28868 2592 28874 2644
rect 32122 2632 32128 2644
rect 32083 2604 32128 2632
rect 32122 2592 32128 2604
rect 32180 2592 32186 2644
rect 58710 2632 58716 2644
rect 32232 2604 58716 2632
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 9732 2536 10241 2564
rect 9732 2524 9738 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 11885 2567 11943 2573
rect 11885 2533 11897 2567
rect 11931 2564 11943 2567
rect 32232 2564 32260 2604
rect 58710 2592 58716 2604
rect 58768 2592 58774 2644
rect 58805 2635 58863 2641
rect 58805 2601 58817 2635
rect 58851 2632 58863 2635
rect 59446 2632 59452 2644
rect 58851 2604 59452 2632
rect 58851 2601 58863 2604
rect 58805 2595 58863 2601
rect 59446 2592 59452 2604
rect 59504 2592 59510 2644
rect 62758 2632 62764 2644
rect 59924 2604 62764 2632
rect 11931 2536 32260 2564
rect 11931 2533 11943 2536
rect 11885 2527 11943 2533
rect 38010 2524 38016 2576
rect 38068 2564 38074 2576
rect 38473 2567 38531 2573
rect 38473 2564 38485 2567
rect 38068 2536 38485 2564
rect 38068 2524 38074 2536
rect 38473 2533 38485 2536
rect 38519 2533 38531 2567
rect 38473 2527 38531 2533
rect 38562 2524 38568 2576
rect 38620 2564 38626 2576
rect 40218 2564 40224 2576
rect 38620 2536 40224 2564
rect 38620 2524 38626 2536
rect 40218 2524 40224 2536
rect 40276 2524 40282 2576
rect 40678 2524 40684 2576
rect 40736 2564 40742 2576
rect 45554 2564 45560 2576
rect 40736 2536 45560 2564
rect 40736 2524 40742 2536
rect 4893 2499 4951 2505
rect 4893 2465 4905 2499
rect 4939 2496 4951 2499
rect 4939 2468 14688 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2682 2428 2688 2440
rect 2643 2400 2688 2428
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 2866 2428 2872 2440
rect 2827 2400 2872 2428
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3292 2400 3985 2428
rect 3292 2388 3298 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 10410 2428 10416 2440
rect 10371 2400 10416 2428
rect 9125 2391 9183 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 12618 2428 12624 2440
rect 12579 2400 12624 2428
rect 11701 2391 11759 2397
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 3053 2363 3111 2369
rect 3053 2329 3065 2363
rect 3099 2360 3111 2363
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 3099 2332 6745 2360
rect 3099 2329 3111 2332
rect 3053 2323 3111 2329
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 6733 2323 6791 2329
rect 10781 2363 10839 2369
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 10962 2360 10968 2372
rect 10827 2332 10968 2360
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 13538 2320 13544 2372
rect 13596 2360 13602 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 13596 2332 14565 2360
rect 13596 2320 13602 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14660 2360 14688 2468
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 27522 2496 27528 2508
rect 16172 2468 27384 2496
rect 27483 2468 27528 2496
rect 16172 2456 16178 2468
rect 15746 2428 15752 2440
rect 15707 2400 15752 2428
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16850 2428 16856 2440
rect 16811 2400 16856 2428
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17460 2400 17693 2428
rect 17460 2388 17466 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2397 18383 2431
rect 19426 2428 19432 2440
rect 19387 2400 19432 2428
rect 18325 2391 18383 2397
rect 18230 2360 18236 2372
rect 14660 2332 18236 2360
rect 14553 2323 14611 2329
rect 18230 2320 18236 2332
rect 18288 2320 18294 2372
rect 18340 2360 18368 2391
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 20036 2400 20085 2428
rect 20036 2388 20042 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 19702 2360 19708 2372
rect 18340 2332 19708 2360
rect 19702 2320 19708 2332
rect 19760 2320 19766 2372
rect 20364 2360 20392 2391
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21968 2400 22201 2428
rect 21968 2388 21974 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 22833 2431 22891 2437
rect 22833 2428 22845 2431
rect 22612 2400 22845 2428
rect 22612 2388 22618 2400
rect 22833 2397 22845 2400
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23477 2431 23535 2437
rect 23477 2428 23489 2431
rect 23256 2400 23489 2428
rect 23256 2388 23262 2400
rect 23477 2397 23489 2400
rect 23523 2397 23535 2431
rect 24670 2428 24676 2440
rect 23477 2391 23535 2397
rect 23584 2400 24676 2428
rect 23584 2360 23612 2400
rect 24670 2388 24676 2400
rect 24728 2388 24734 2440
rect 24765 2431 24823 2437
rect 24765 2397 24777 2431
rect 24811 2428 24823 2431
rect 24854 2428 24860 2440
rect 24811 2400 24860 2428
rect 24811 2397 24823 2400
rect 24765 2391 24823 2397
rect 24854 2388 24860 2400
rect 24912 2388 24918 2440
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 25188 2400 25237 2428
rect 25188 2388 25194 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2428 26479 2431
rect 27062 2428 27068 2440
rect 26467 2400 27068 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 27062 2388 27068 2400
rect 27120 2388 27126 2440
rect 27356 2437 27384 2468
rect 27522 2456 27528 2468
rect 27580 2456 27586 2508
rect 29730 2496 29736 2508
rect 27816 2468 29736 2496
rect 27341 2431 27399 2437
rect 27341 2397 27353 2431
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 27433 2431 27491 2437
rect 27433 2397 27445 2431
rect 27479 2424 27491 2431
rect 27706 2428 27712 2440
rect 27540 2424 27712 2428
rect 27479 2400 27712 2424
rect 27479 2397 27568 2400
rect 27433 2396 27568 2397
rect 27433 2391 27491 2396
rect 27706 2388 27712 2400
rect 27764 2388 27770 2440
rect 27816 2360 27844 2468
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 29822 2456 29828 2508
rect 29880 2496 29886 2508
rect 32766 2496 32772 2508
rect 29880 2468 32628 2496
rect 32727 2468 32772 2496
rect 29880 2456 29886 2468
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 28810 2428 28816 2440
rect 28399 2400 28816 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 28810 2388 28816 2400
rect 28868 2388 28874 2440
rect 28994 2428 29000 2440
rect 28955 2400 29000 2428
rect 28994 2388 29000 2400
rect 29052 2388 29058 2440
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29696 2400 29929 2428
rect 29696 2388 29702 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 30926 2428 30932 2440
rect 30887 2400 30932 2428
rect 29917 2391 29975 2397
rect 30926 2388 30932 2400
rect 30984 2388 30990 2440
rect 31570 2428 31576 2440
rect 31531 2400 31576 2428
rect 31570 2388 31576 2400
rect 31628 2388 31634 2440
rect 20364 2332 23612 2360
rect 27356 2332 27844 2360
rect 27356 2304 27384 2332
rect 28258 2320 28264 2372
rect 28316 2360 28322 2372
rect 32600 2369 32628 2468
rect 32766 2456 32772 2468
rect 32824 2456 32830 2508
rect 34698 2496 34704 2508
rect 33336 2468 33916 2496
rect 34659 2468 34704 2496
rect 32493 2363 32551 2369
rect 32493 2360 32505 2363
rect 28316 2332 32505 2360
rect 28316 2320 28322 2332
rect 32493 2329 32505 2332
rect 32539 2329 32551 2363
rect 32493 2323 32551 2329
rect 32585 2363 32643 2369
rect 32585 2329 32597 2363
rect 32631 2360 32643 2363
rect 33137 2363 33195 2369
rect 33137 2360 33149 2363
rect 32631 2332 33149 2360
rect 32631 2329 32643 2332
rect 32585 2323 32643 2329
rect 33137 2329 33149 2332
rect 33183 2329 33195 2363
rect 33137 2323 33195 2329
rect 7006 2292 7012 2304
rect 6967 2264 7012 2292
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 8205 2295 8263 2301
rect 8205 2261 8217 2295
rect 8251 2292 8263 2295
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 8251 2264 8585 2292
rect 8251 2261 8263 2264
rect 8205 2255 8263 2261
rect 8573 2261 8585 2264
rect 8619 2292 8631 2295
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 8619 2264 9321 2292
rect 8619 2261 8631 2264
rect 8573 2255 8631 2261
rect 9309 2261 9321 2264
rect 9355 2292 9367 2295
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9355 2264 9781 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 9769 2261 9781 2264
rect 9815 2292 9827 2295
rect 10134 2292 10140 2304
rect 9815 2264 10140 2292
rect 9815 2261 9827 2264
rect 9769 2255 9827 2261
rect 10134 2252 10140 2264
rect 10192 2252 10198 2304
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12308 2264 12449 2292
rect 12308 2252 12314 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15565 2295 15623 2301
rect 15565 2292 15577 2295
rect 15528 2264 15577 2292
rect 15528 2252 15534 2264
rect 15565 2261 15577 2264
rect 15611 2261 15623 2295
rect 15565 2255 15623 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16669 2295 16727 2301
rect 16669 2292 16681 2295
rect 16172 2264 16681 2292
rect 16172 2252 16178 2264
rect 16669 2261 16681 2264
rect 16715 2261 16727 2295
rect 17494 2292 17500 2304
rect 17455 2264 17500 2292
rect 16669 2255 16727 2261
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18141 2295 18199 2301
rect 18141 2292 18153 2295
rect 18104 2264 18153 2292
rect 18104 2252 18110 2264
rect 18141 2261 18153 2264
rect 18187 2261 18199 2295
rect 18141 2255 18199 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 19245 2295 19303 2301
rect 19245 2292 19257 2295
rect 18748 2264 19257 2292
rect 18748 2252 18754 2264
rect 19245 2261 19257 2264
rect 19291 2261 19303 2295
rect 19245 2255 19303 2261
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24544 2264 24593 2292
rect 24544 2252 24550 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 24670 2252 24676 2304
rect 24728 2292 24734 2304
rect 26142 2292 26148 2304
rect 24728 2264 26148 2292
rect 24728 2252 24734 2264
rect 26142 2252 26148 2264
rect 26200 2252 26206 2304
rect 26237 2295 26295 2301
rect 26237 2261 26249 2295
rect 26283 2292 26295 2295
rect 27154 2292 27160 2304
rect 26283 2264 27160 2292
rect 26283 2261 26295 2264
rect 26237 2255 26295 2261
rect 27154 2252 27160 2264
rect 27212 2252 27218 2304
rect 27338 2252 27344 2304
rect 27396 2252 27402 2304
rect 28166 2292 28172 2304
rect 28127 2264 28172 2292
rect 28166 2252 28172 2264
rect 28224 2252 28230 2304
rect 29730 2292 29736 2304
rect 29691 2264 29736 2292
rect 29730 2252 29736 2264
rect 29788 2252 29794 2304
rect 30742 2292 30748 2304
rect 30703 2264 30748 2292
rect 30742 2252 30748 2264
rect 30800 2252 30806 2304
rect 31294 2252 31300 2304
rect 31352 2292 31358 2304
rect 31389 2295 31447 2301
rect 31389 2292 31401 2295
rect 31352 2264 31401 2292
rect 31352 2252 31358 2264
rect 31389 2261 31401 2264
rect 31435 2261 31447 2295
rect 31389 2255 31447 2261
rect 31662 2252 31668 2304
rect 31720 2292 31726 2304
rect 33336 2292 33364 2468
rect 33781 2431 33839 2437
rect 33781 2397 33793 2431
rect 33827 2397 33839 2431
rect 33888 2428 33916 2468
rect 34698 2456 34704 2468
rect 34756 2456 34762 2508
rect 36633 2499 36691 2505
rect 36633 2465 36645 2499
rect 36679 2496 36691 2499
rect 37826 2496 37832 2508
rect 36679 2468 37832 2496
rect 36679 2465 36691 2468
rect 36633 2459 36691 2465
rect 37826 2456 37832 2468
rect 37884 2456 37890 2508
rect 40788 2505 40816 2536
rect 45554 2524 45560 2536
rect 45612 2524 45618 2576
rect 47578 2564 47584 2576
rect 47539 2536 47584 2564
rect 47578 2524 47584 2536
rect 47636 2524 47642 2576
rect 50430 2564 50436 2576
rect 47872 2536 50436 2564
rect 40773 2499 40831 2505
rect 40773 2465 40785 2499
rect 40819 2465 40831 2499
rect 40773 2459 40831 2465
rect 42429 2499 42487 2505
rect 42429 2465 42441 2499
rect 42475 2496 42487 2499
rect 42610 2496 42616 2508
rect 42475 2468 42616 2496
rect 42475 2465 42487 2468
rect 42429 2459 42487 2465
rect 42610 2456 42616 2468
rect 42668 2456 42674 2508
rect 46750 2496 46756 2508
rect 46711 2468 46756 2496
rect 46750 2456 46756 2468
rect 46808 2456 46814 2508
rect 46937 2499 46995 2505
rect 46937 2465 46949 2499
rect 46983 2496 46995 2499
rect 47872 2496 47900 2536
rect 48038 2496 48044 2508
rect 46983 2468 47900 2496
rect 47999 2468 48044 2496
rect 46983 2465 46995 2468
rect 46937 2459 46995 2465
rect 48038 2456 48044 2468
rect 48096 2456 48102 2508
rect 48240 2505 48268 2536
rect 50430 2524 50436 2536
rect 50488 2524 50494 2576
rect 50798 2524 50804 2576
rect 50856 2564 50862 2576
rect 52730 2564 52736 2576
rect 50856 2536 52132 2564
rect 52691 2536 52736 2564
rect 50856 2524 50862 2536
rect 48225 2499 48283 2505
rect 48225 2465 48237 2499
rect 48271 2465 48283 2499
rect 51994 2496 52000 2508
rect 48225 2459 48283 2465
rect 50356 2468 51764 2496
rect 51955 2468 52000 2496
rect 34977 2431 35035 2437
rect 34977 2428 34989 2431
rect 33888 2400 34989 2428
rect 33781 2391 33839 2397
rect 34977 2397 34989 2400
rect 35023 2397 35035 2431
rect 34977 2391 35035 2397
rect 35912 2400 36216 2428
rect 33796 2360 33824 2391
rect 35912 2360 35940 2400
rect 33796 2332 35940 2360
rect 31720 2264 33364 2292
rect 31720 2252 31726 2264
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33597 2295 33655 2301
rect 33597 2292 33609 2295
rect 33560 2264 33609 2292
rect 33560 2252 33566 2264
rect 33597 2261 33609 2264
rect 33643 2261 33655 2295
rect 33597 2255 33655 2261
rect 34698 2252 34704 2304
rect 34756 2292 34762 2304
rect 35989 2295 36047 2301
rect 35989 2292 36001 2295
rect 34756 2264 36001 2292
rect 34756 2252 34762 2264
rect 35989 2261 36001 2264
rect 36035 2261 36047 2295
rect 36188 2292 36216 2400
rect 36262 2388 36268 2440
rect 36320 2428 36326 2440
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 36320 2400 36369 2428
rect 36320 2388 36326 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 37642 2428 37648 2440
rect 37603 2400 37648 2428
rect 36357 2391 36415 2397
rect 37642 2388 37648 2400
rect 37700 2388 37706 2440
rect 38197 2431 38255 2437
rect 38197 2397 38209 2431
rect 38243 2428 38255 2431
rect 38654 2428 38660 2440
rect 38243 2400 38660 2428
rect 38243 2397 38255 2400
rect 38197 2391 38255 2397
rect 38654 2388 38660 2400
rect 38712 2388 38718 2440
rect 39298 2428 39304 2440
rect 39259 2400 39304 2428
rect 39298 2388 39304 2400
rect 39356 2388 39362 2440
rect 40126 2388 40132 2440
rect 40184 2428 40190 2440
rect 40497 2431 40555 2437
rect 40497 2428 40509 2431
rect 40184 2400 40509 2428
rect 40184 2388 40190 2400
rect 40497 2397 40509 2400
rect 40543 2397 40555 2431
rect 42702 2428 42708 2440
rect 42663 2400 42708 2428
rect 40497 2391 40555 2397
rect 42702 2388 42708 2400
rect 42760 2388 42766 2440
rect 44453 2431 44511 2437
rect 44453 2397 44465 2431
rect 44499 2428 44511 2431
rect 45922 2428 45928 2440
rect 44499 2400 45928 2428
rect 44499 2397 44511 2400
rect 44453 2391 44511 2397
rect 45922 2388 45928 2400
rect 45980 2388 45986 2440
rect 46017 2431 46075 2437
rect 46017 2397 46029 2431
rect 46063 2428 46075 2431
rect 46063 2400 46704 2428
rect 46063 2397 46075 2400
rect 46017 2391 46075 2397
rect 36449 2363 36507 2369
rect 36449 2329 36461 2363
rect 36495 2360 36507 2363
rect 36538 2360 36544 2372
rect 36495 2332 36544 2360
rect 36495 2329 36507 2332
rect 36449 2323 36507 2329
rect 36538 2320 36544 2332
rect 36596 2320 36602 2372
rect 39850 2360 39856 2372
rect 37292 2332 39856 2360
rect 37292 2292 37320 2332
rect 39850 2320 39856 2332
rect 39908 2320 39914 2372
rect 41601 2363 41659 2369
rect 41601 2360 41613 2363
rect 40144 2332 41613 2360
rect 36188 2264 37320 2292
rect 35989 2255 36047 2261
rect 37366 2252 37372 2304
rect 37424 2292 37430 2304
rect 37461 2295 37519 2301
rect 37461 2292 37473 2295
rect 37424 2264 37473 2292
rect 37424 2252 37430 2264
rect 37461 2261 37473 2264
rect 37507 2261 37519 2295
rect 37461 2255 37519 2261
rect 39117 2295 39175 2301
rect 39117 2261 39129 2295
rect 39163 2292 39175 2295
rect 39942 2292 39948 2304
rect 39163 2264 39948 2292
rect 39163 2261 39175 2264
rect 39117 2255 39175 2261
rect 39942 2252 39948 2264
rect 40000 2252 40006 2304
rect 40144 2301 40172 2332
rect 41601 2329 41613 2332
rect 41647 2329 41659 2363
rect 41782 2360 41788 2372
rect 41743 2332 41788 2360
rect 41601 2323 41659 2329
rect 41782 2320 41788 2332
rect 41840 2320 41846 2372
rect 45465 2363 45523 2369
rect 45465 2329 45477 2363
rect 45511 2360 45523 2363
rect 45511 2332 46336 2360
rect 45511 2329 45523 2332
rect 45465 2323 45523 2329
rect 40129 2295 40187 2301
rect 40129 2261 40141 2295
rect 40175 2261 40187 2295
rect 40129 2255 40187 2261
rect 40494 2252 40500 2304
rect 40552 2292 40558 2304
rect 40589 2295 40647 2301
rect 40589 2292 40601 2295
rect 40552 2264 40601 2292
rect 40552 2252 40558 2264
rect 40589 2261 40601 2264
rect 40635 2292 40647 2295
rect 41141 2295 41199 2301
rect 41141 2292 41153 2295
rect 40635 2264 41153 2292
rect 40635 2261 40647 2264
rect 40589 2255 40647 2261
rect 41141 2261 41153 2264
rect 41187 2261 41199 2295
rect 41141 2255 41199 2261
rect 44269 2295 44327 2301
rect 44269 2261 44281 2295
rect 44315 2292 44327 2295
rect 44450 2292 44456 2304
rect 44315 2264 44456 2292
rect 44315 2261 44327 2264
rect 44269 2255 44327 2261
rect 44450 2252 44456 2264
rect 44508 2252 44514 2304
rect 45554 2252 45560 2304
rect 45612 2292 45618 2304
rect 46308 2301 46336 2332
rect 46676 2304 46704 2400
rect 49142 2388 49148 2440
rect 49200 2428 49206 2440
rect 50356 2437 50384 2468
rect 49237 2431 49295 2437
rect 49237 2428 49249 2431
rect 49200 2400 49249 2428
rect 49200 2388 49206 2400
rect 49237 2397 49249 2400
rect 49283 2397 49295 2431
rect 49237 2391 49295 2397
rect 50341 2431 50399 2437
rect 50341 2397 50353 2431
rect 50387 2397 50399 2431
rect 50341 2391 50399 2397
rect 50985 2431 51043 2437
rect 50985 2397 50997 2431
rect 51031 2428 51043 2431
rect 51736 2428 51764 2468
rect 51994 2456 52000 2468
rect 52052 2456 52058 2508
rect 52104 2496 52132 2536
rect 52730 2524 52736 2536
rect 52788 2524 52794 2576
rect 54018 2564 54024 2576
rect 52840 2536 54024 2564
rect 52840 2496 52868 2536
rect 52104 2468 52868 2496
rect 52914 2456 52920 2508
rect 52972 2496 52978 2508
rect 53300 2505 53328 2536
rect 54018 2524 54024 2536
rect 54076 2524 54082 2576
rect 54573 2567 54631 2573
rect 54573 2533 54585 2567
rect 54619 2564 54631 2567
rect 59924 2564 59952 2604
rect 62758 2592 62764 2604
rect 62816 2592 62822 2644
rect 63770 2592 63776 2644
rect 63828 2632 63834 2644
rect 64509 2635 64567 2641
rect 64509 2632 64521 2635
rect 63828 2604 64521 2632
rect 63828 2592 63834 2604
rect 64509 2601 64521 2604
rect 64555 2601 64567 2635
rect 66714 2632 66720 2644
rect 66675 2604 66720 2632
rect 64509 2595 64567 2601
rect 66714 2592 66720 2604
rect 66772 2592 66778 2644
rect 70762 2632 70768 2644
rect 66824 2604 70624 2632
rect 70723 2604 70768 2632
rect 54619 2536 59952 2564
rect 54619 2533 54631 2536
rect 54573 2527 54631 2533
rect 59998 2524 60004 2576
rect 60056 2564 60062 2576
rect 60645 2567 60703 2573
rect 60645 2564 60657 2567
rect 60056 2536 60657 2564
rect 60056 2524 60062 2536
rect 60645 2533 60657 2536
rect 60691 2533 60703 2567
rect 60645 2527 60703 2533
rect 61120 2536 61516 2564
rect 53193 2499 53251 2505
rect 53193 2496 53205 2499
rect 52972 2468 53205 2496
rect 52972 2456 52978 2468
rect 53193 2465 53205 2468
rect 53239 2465 53251 2499
rect 53193 2459 53251 2465
rect 53285 2499 53343 2505
rect 53285 2465 53297 2499
rect 53331 2465 53343 2499
rect 56410 2496 56416 2508
rect 53285 2459 53343 2465
rect 53392 2468 56416 2496
rect 53392 2428 53420 2468
rect 56410 2456 56416 2468
rect 56468 2456 56474 2508
rect 56778 2496 56784 2508
rect 56739 2468 56784 2496
rect 56778 2456 56784 2468
rect 56836 2456 56842 2508
rect 57790 2456 57796 2508
rect 57848 2496 57854 2508
rect 59265 2499 59323 2505
rect 59265 2496 59277 2499
rect 57848 2468 59277 2496
rect 57848 2456 57854 2468
rect 59265 2465 59277 2468
rect 59311 2465 59323 2499
rect 59265 2459 59323 2465
rect 59449 2499 59507 2505
rect 59449 2465 59461 2499
rect 59495 2496 59507 2499
rect 61120 2496 61148 2536
rect 59495 2468 61148 2496
rect 61197 2499 61255 2505
rect 59495 2465 59507 2468
rect 59449 2459 59507 2465
rect 61197 2465 61209 2499
rect 61243 2496 61255 2499
rect 61488 2496 61516 2536
rect 62574 2524 62580 2576
rect 62632 2564 62638 2576
rect 66824 2564 66852 2604
rect 62632 2536 66852 2564
rect 66916 2536 67404 2564
rect 62632 2524 62638 2536
rect 66916 2496 66944 2536
rect 67269 2499 67327 2505
rect 67269 2496 67281 2499
rect 61243 2468 61332 2496
rect 61488 2468 66944 2496
rect 67008 2468 67281 2496
rect 61243 2465 61255 2468
rect 61197 2459 61255 2465
rect 51031 2400 51488 2428
rect 51736 2400 53420 2428
rect 51031 2397 51043 2400
rect 50985 2391 51043 2397
rect 46750 2320 46756 2372
rect 46808 2360 46814 2372
rect 46808 2332 50844 2360
rect 46808 2320 46814 2332
rect 46293 2295 46351 2301
rect 45612 2264 45657 2292
rect 45612 2252 45618 2264
rect 46293 2261 46305 2295
rect 46339 2261 46351 2295
rect 46658 2292 46664 2304
rect 46619 2264 46664 2292
rect 46293 2255 46351 2261
rect 46658 2252 46664 2264
rect 46716 2252 46722 2304
rect 47946 2292 47952 2304
rect 47907 2264 47952 2292
rect 47946 2252 47952 2264
rect 48004 2252 48010 2304
rect 48958 2252 48964 2304
rect 49016 2292 49022 2304
rect 49053 2295 49111 2301
rect 49053 2292 49065 2295
rect 49016 2264 49065 2292
rect 49016 2252 49022 2264
rect 49053 2261 49065 2264
rect 49099 2261 49111 2295
rect 49053 2255 49111 2261
rect 50157 2295 50215 2301
rect 50157 2261 50169 2295
rect 50203 2292 50215 2295
rect 50246 2292 50252 2304
rect 50203 2264 50252 2292
rect 50203 2261 50215 2264
rect 50157 2255 50215 2261
rect 50246 2252 50252 2264
rect 50304 2252 50310 2304
rect 50816 2301 50844 2332
rect 51460 2301 51488 2400
rect 53926 2388 53932 2440
rect 53984 2388 53990 2440
rect 54110 2428 54116 2440
rect 54071 2400 54116 2428
rect 54110 2388 54116 2400
rect 54168 2388 54174 2440
rect 54754 2428 54760 2440
rect 54715 2400 54760 2428
rect 54754 2388 54760 2400
rect 54812 2388 54818 2440
rect 56505 2431 56563 2437
rect 55186 2400 55996 2428
rect 51626 2320 51632 2372
rect 51684 2360 51690 2372
rect 53944 2360 53972 2388
rect 51684 2332 53972 2360
rect 51684 2320 51690 2332
rect 54018 2320 54024 2372
rect 54076 2360 54082 2372
rect 55186 2360 55214 2400
rect 55858 2360 55864 2372
rect 54076 2332 55214 2360
rect 55819 2332 55864 2360
rect 54076 2320 54082 2332
rect 55858 2320 55864 2332
rect 55916 2320 55922 2372
rect 55968 2360 55996 2400
rect 56505 2397 56517 2431
rect 56551 2428 56563 2431
rect 56686 2428 56692 2440
rect 56551 2400 56692 2428
rect 56551 2397 56563 2400
rect 56505 2391 56563 2397
rect 56686 2388 56692 2400
rect 56744 2388 56750 2440
rect 58158 2428 58164 2440
rect 58119 2400 58164 2428
rect 58158 2388 58164 2400
rect 58216 2388 58222 2440
rect 59464 2428 59492 2459
rect 61304 2440 61332 2468
rect 59096 2400 59492 2428
rect 59096 2360 59124 2400
rect 61286 2388 61292 2440
rect 61344 2388 61350 2440
rect 61470 2388 61476 2440
rect 61528 2428 61534 2440
rect 62025 2431 62083 2437
rect 62025 2428 62037 2431
rect 61528 2400 62037 2428
rect 61528 2388 61534 2400
rect 62025 2397 62037 2400
rect 62071 2397 62083 2431
rect 63402 2428 63408 2440
rect 63363 2400 63408 2428
rect 62025 2391 62083 2397
rect 63402 2388 63408 2400
rect 63460 2388 63466 2440
rect 64046 2428 64052 2440
rect 64007 2400 64052 2428
rect 64046 2388 64052 2400
rect 64104 2388 64110 2440
rect 64693 2431 64751 2437
rect 64693 2397 64705 2431
rect 64739 2397 64751 2431
rect 65978 2428 65984 2440
rect 65939 2400 65984 2428
rect 64693 2391 64751 2397
rect 55968 2332 59124 2360
rect 59173 2363 59231 2369
rect 59173 2329 59185 2363
rect 59219 2360 59231 2363
rect 59354 2360 59360 2372
rect 59219 2332 59360 2360
rect 59219 2329 59231 2332
rect 59173 2323 59231 2329
rect 59354 2320 59360 2332
rect 59412 2320 59418 2372
rect 64708 2360 64736 2391
rect 65978 2388 65984 2400
rect 66036 2388 66042 2440
rect 66070 2388 66076 2440
rect 66128 2428 66134 2440
rect 67008 2428 67036 2468
rect 67269 2465 67281 2468
rect 67315 2465 67327 2499
rect 67376 2496 67404 2536
rect 67450 2524 67456 2576
rect 67508 2564 67514 2576
rect 68557 2567 68615 2573
rect 68557 2564 68569 2567
rect 67508 2536 68569 2564
rect 67508 2524 67514 2536
rect 68557 2533 68569 2536
rect 68603 2564 68615 2567
rect 68922 2564 68928 2576
rect 68603 2536 68928 2564
rect 68603 2533 68615 2536
rect 68557 2527 68615 2533
rect 68922 2524 68928 2536
rect 68980 2524 68986 2576
rect 69293 2567 69351 2573
rect 69293 2533 69305 2567
rect 69339 2564 69351 2567
rect 70394 2564 70400 2576
rect 69339 2536 70400 2564
rect 69339 2533 69351 2536
rect 69293 2527 69351 2533
rect 70394 2524 70400 2536
rect 70452 2524 70458 2576
rect 70596 2564 70624 2604
rect 70762 2592 70768 2604
rect 70820 2592 70826 2644
rect 71314 2592 71320 2644
rect 71372 2632 71378 2644
rect 71593 2635 71651 2641
rect 71593 2632 71605 2635
rect 71372 2604 71605 2632
rect 71372 2592 71378 2604
rect 71593 2601 71605 2604
rect 71639 2601 71651 2635
rect 71593 2595 71651 2601
rect 72326 2592 72332 2644
rect 72384 2632 72390 2644
rect 72605 2635 72663 2641
rect 72605 2632 72617 2635
rect 72384 2604 72617 2632
rect 72384 2592 72390 2604
rect 72605 2601 72617 2604
rect 72651 2601 72663 2635
rect 82446 2632 82452 2644
rect 72605 2595 72663 2601
rect 73816 2604 82452 2632
rect 73816 2564 73844 2604
rect 82446 2592 82452 2604
rect 82504 2592 82510 2644
rect 82538 2592 82544 2644
rect 82596 2632 82602 2644
rect 82596 2604 82641 2632
rect 82596 2592 82602 2604
rect 82722 2592 82728 2644
rect 82780 2632 82786 2644
rect 100205 2635 100263 2641
rect 100205 2632 100217 2635
rect 82780 2604 100217 2632
rect 82780 2592 82786 2604
rect 100205 2601 100217 2604
rect 100251 2632 100263 2635
rect 100757 2635 100815 2641
rect 100757 2632 100769 2635
rect 100251 2604 100769 2632
rect 100251 2601 100263 2604
rect 100205 2595 100263 2601
rect 100757 2601 100769 2604
rect 100803 2601 100815 2635
rect 102226 2632 102232 2644
rect 102187 2604 102232 2632
rect 100757 2595 100815 2601
rect 102226 2592 102232 2604
rect 102284 2592 102290 2644
rect 103330 2632 103336 2644
rect 103291 2604 103336 2632
rect 103330 2592 103336 2604
rect 103388 2592 103394 2644
rect 104526 2592 104532 2644
rect 104584 2632 104590 2644
rect 111061 2635 111119 2641
rect 111061 2632 111073 2635
rect 104584 2604 111073 2632
rect 104584 2592 104590 2604
rect 111061 2601 111073 2604
rect 111107 2601 111119 2635
rect 111061 2595 111119 2601
rect 114557 2635 114615 2641
rect 114557 2601 114569 2635
rect 114603 2632 114615 2635
rect 114738 2632 114744 2644
rect 114603 2604 114744 2632
rect 114603 2601 114615 2604
rect 114557 2595 114615 2601
rect 114738 2592 114744 2604
rect 114796 2592 114802 2644
rect 118234 2564 118240 2576
rect 70596 2536 73844 2564
rect 73908 2536 82492 2564
rect 69845 2499 69903 2505
rect 69845 2496 69857 2499
rect 67376 2468 69857 2496
rect 67269 2459 67327 2465
rect 69845 2465 69857 2468
rect 69891 2465 69903 2499
rect 69845 2459 69903 2465
rect 66128 2400 67036 2428
rect 66128 2388 66134 2400
rect 67358 2388 67364 2440
rect 67416 2428 67422 2440
rect 68005 2431 68063 2437
rect 68005 2428 68017 2431
rect 67416 2424 67496 2428
rect 67560 2424 68017 2428
rect 67416 2400 68017 2424
rect 67416 2388 67422 2400
rect 67468 2396 67588 2400
rect 68005 2397 68017 2400
rect 68051 2397 68063 2431
rect 69658 2428 69664 2440
rect 69619 2400 69664 2428
rect 68005 2391 68063 2397
rect 69658 2388 69664 2400
rect 69716 2388 69722 2440
rect 69860 2428 69888 2459
rect 69934 2456 69940 2508
rect 69992 2496 69998 2508
rect 71866 2496 71872 2508
rect 69992 2468 71872 2496
rect 69992 2456 69998 2468
rect 71866 2456 71872 2468
rect 71924 2456 71930 2508
rect 72050 2496 72056 2508
rect 72011 2468 72056 2496
rect 72050 2456 72056 2468
rect 72108 2456 72114 2508
rect 72145 2499 72203 2505
rect 72145 2465 72157 2499
rect 72191 2465 72203 2499
rect 72145 2459 72203 2465
rect 70578 2428 70584 2440
rect 69860 2400 70584 2428
rect 70578 2388 70584 2400
rect 70636 2388 70642 2440
rect 70949 2431 71007 2437
rect 70949 2397 70961 2431
rect 70995 2428 71007 2431
rect 71222 2428 71228 2440
rect 70995 2400 71228 2428
rect 70995 2397 71007 2400
rect 70949 2391 71007 2397
rect 71222 2388 71228 2400
rect 71280 2388 71286 2440
rect 71314 2388 71320 2440
rect 71372 2428 71378 2440
rect 72160 2428 72188 2459
rect 73522 2456 73528 2508
rect 73580 2496 73586 2508
rect 73908 2496 73936 2536
rect 73580 2468 73936 2496
rect 73580 2456 73586 2468
rect 73982 2456 73988 2508
rect 74040 2496 74046 2508
rect 74040 2468 74085 2496
rect 74040 2456 74046 2468
rect 77018 2456 77024 2508
rect 77076 2496 77082 2508
rect 77113 2499 77171 2505
rect 77113 2496 77125 2499
rect 77076 2468 77125 2496
rect 77076 2456 77082 2468
rect 77113 2465 77125 2468
rect 77159 2465 77171 2499
rect 77113 2459 77171 2465
rect 77202 2456 77208 2508
rect 77260 2496 77266 2508
rect 82464 2496 82492 2536
rect 82648 2536 118240 2564
rect 82648 2496 82676 2536
rect 118234 2524 118240 2536
rect 118292 2524 118298 2576
rect 77260 2468 81572 2496
rect 82464 2468 82676 2496
rect 77260 2456 77266 2468
rect 71372 2400 72188 2428
rect 71372 2388 71378 2400
rect 73706 2388 73712 2440
rect 73764 2428 73770 2440
rect 73803 2431 73861 2437
rect 73803 2428 73815 2431
rect 73764 2400 73815 2428
rect 73764 2388 73770 2400
rect 73803 2397 73815 2400
rect 73849 2397 73861 2431
rect 73803 2391 73861 2397
rect 74445 2431 74503 2437
rect 74445 2397 74457 2431
rect 74491 2428 74503 2431
rect 75733 2431 75791 2437
rect 74491 2400 75684 2428
rect 74491 2397 74503 2400
rect 74445 2391 74503 2397
rect 63880 2332 64736 2360
rect 50801 2295 50859 2301
rect 50801 2261 50813 2295
rect 50847 2261 50859 2295
rect 50801 2255 50859 2261
rect 51445 2295 51503 2301
rect 51445 2261 51457 2295
rect 51491 2261 51503 2295
rect 51810 2292 51816 2304
rect 51771 2264 51816 2292
rect 51445 2255 51503 2261
rect 51810 2252 51816 2264
rect 51868 2252 51874 2304
rect 51902 2252 51908 2304
rect 51960 2292 51966 2304
rect 53098 2292 53104 2304
rect 51960 2264 52005 2292
rect 53059 2264 53104 2292
rect 51960 2252 51966 2264
rect 53098 2252 53104 2264
rect 53156 2252 53162 2304
rect 53466 2252 53472 2304
rect 53524 2292 53530 2304
rect 53929 2295 53987 2301
rect 53929 2292 53941 2295
rect 53524 2264 53941 2292
rect 53524 2252 53530 2264
rect 53929 2261 53941 2264
rect 53975 2261 53987 2295
rect 55950 2292 55956 2304
rect 55911 2264 55956 2292
rect 53929 2255 53987 2261
rect 55950 2252 55956 2264
rect 56008 2252 56014 2304
rect 58250 2292 58256 2304
rect 58211 2264 58256 2292
rect 58250 2252 58256 2264
rect 58308 2252 58314 2304
rect 61010 2292 61016 2304
rect 60971 2264 61016 2292
rect 61010 2252 61016 2264
rect 61068 2252 61074 2304
rect 61105 2295 61163 2301
rect 61105 2261 61117 2295
rect 61151 2292 61163 2295
rect 61841 2295 61899 2301
rect 61841 2292 61853 2295
rect 61151 2264 61853 2292
rect 61151 2261 61163 2264
rect 61105 2255 61163 2261
rect 61841 2261 61853 2264
rect 61887 2261 61899 2295
rect 61841 2255 61899 2261
rect 63126 2252 63132 2304
rect 63184 2292 63190 2304
rect 63880 2301 63908 2332
rect 66806 2320 66812 2372
rect 66864 2360 66870 2372
rect 67085 2363 67143 2369
rect 67085 2360 67097 2363
rect 66864 2332 67097 2360
rect 66864 2320 66870 2332
rect 67085 2329 67097 2332
rect 67131 2329 67143 2363
rect 67085 2323 67143 2329
rect 67266 2320 67272 2372
rect 67324 2360 67330 2372
rect 71038 2360 71044 2372
rect 67324 2332 71044 2360
rect 67324 2320 67330 2332
rect 71038 2320 71044 2332
rect 71096 2320 71102 2372
rect 71130 2320 71136 2372
rect 71188 2360 71194 2372
rect 71188 2332 73752 2360
rect 71188 2320 71194 2332
rect 63221 2295 63279 2301
rect 63221 2292 63233 2295
rect 63184 2264 63233 2292
rect 63184 2252 63190 2264
rect 63221 2261 63233 2264
rect 63267 2261 63279 2295
rect 63221 2255 63279 2261
rect 63865 2295 63923 2301
rect 63865 2261 63877 2295
rect 63911 2261 63923 2295
rect 63865 2255 63923 2261
rect 65702 2252 65708 2304
rect 65760 2292 65766 2304
rect 65797 2295 65855 2301
rect 65797 2292 65809 2295
rect 65760 2264 65809 2292
rect 65760 2252 65766 2264
rect 65797 2261 65809 2264
rect 65843 2261 65855 2295
rect 65797 2255 65855 2261
rect 66441 2295 66499 2301
rect 66441 2261 66453 2295
rect 66487 2292 66499 2295
rect 67174 2292 67180 2304
rect 66487 2264 67180 2292
rect 66487 2261 66499 2264
rect 66441 2255 66499 2261
rect 67174 2252 67180 2264
rect 67232 2292 67238 2304
rect 67232 2264 67325 2292
rect 67232 2252 67238 2264
rect 67634 2252 67640 2304
rect 67692 2292 67698 2304
rect 67821 2295 67879 2301
rect 67821 2292 67833 2295
rect 67692 2264 67833 2292
rect 67692 2252 67698 2264
rect 67821 2261 67833 2264
rect 67867 2261 67879 2295
rect 67821 2255 67879 2261
rect 68922 2252 68928 2304
rect 68980 2292 68986 2304
rect 69753 2295 69811 2301
rect 69753 2292 69765 2295
rect 68980 2264 69765 2292
rect 68980 2252 68986 2264
rect 69753 2261 69765 2264
rect 69799 2292 69811 2295
rect 70305 2295 70363 2301
rect 70305 2292 70317 2295
rect 69799 2264 70317 2292
rect 69799 2261 69811 2264
rect 69753 2255 69811 2261
rect 70305 2261 70317 2264
rect 70351 2292 70363 2295
rect 71225 2295 71283 2301
rect 71225 2292 71237 2295
rect 70351 2264 71237 2292
rect 70351 2261 70363 2264
rect 70305 2255 70363 2261
rect 71225 2261 71237 2264
rect 71271 2261 71283 2295
rect 71225 2255 71283 2261
rect 71961 2295 72019 2301
rect 71961 2261 71973 2295
rect 72007 2292 72019 2295
rect 73614 2292 73620 2304
rect 72007 2264 73620 2292
rect 72007 2261 72019 2264
rect 71961 2255 72019 2261
rect 73614 2252 73620 2264
rect 73672 2252 73678 2304
rect 73724 2292 73752 2332
rect 73908 2332 75592 2360
rect 73908 2292 73936 2332
rect 74626 2292 74632 2304
rect 73724 2264 73936 2292
rect 74587 2264 74632 2292
rect 74626 2252 74632 2264
rect 74684 2252 74690 2304
rect 75564 2301 75592 2332
rect 75549 2295 75607 2301
rect 75549 2261 75561 2295
rect 75595 2261 75607 2295
rect 75656 2292 75684 2400
rect 75733 2397 75745 2431
rect 75779 2428 75791 2431
rect 75822 2428 75828 2440
rect 75779 2400 75828 2428
rect 75779 2397 75791 2400
rect 75733 2391 75791 2397
rect 75822 2388 75828 2400
rect 75880 2388 75886 2440
rect 77386 2388 77392 2440
rect 77444 2428 77450 2440
rect 77941 2431 77999 2437
rect 77941 2428 77953 2431
rect 77444 2400 77953 2428
rect 77444 2388 77450 2400
rect 77941 2397 77953 2400
rect 77987 2397 77999 2431
rect 77941 2391 77999 2397
rect 78030 2388 78036 2440
rect 78088 2428 78094 2440
rect 78861 2431 78919 2437
rect 78861 2428 78873 2431
rect 78088 2400 78873 2428
rect 78088 2388 78094 2400
rect 78861 2397 78873 2400
rect 78907 2397 78919 2431
rect 79502 2428 79508 2440
rect 79463 2400 79508 2428
rect 78861 2391 78919 2397
rect 79502 2388 79508 2400
rect 79560 2388 79566 2440
rect 80514 2388 80520 2440
rect 80572 2428 80578 2440
rect 81069 2431 81127 2437
rect 81069 2428 81081 2431
rect 80572 2400 81081 2428
rect 80572 2388 80578 2400
rect 81069 2397 81081 2400
rect 81115 2397 81127 2431
rect 81342 2428 81348 2440
rect 81303 2400 81348 2428
rect 81069 2391 81127 2397
rect 81342 2388 81348 2400
rect 81400 2388 81406 2440
rect 81544 2428 81572 2468
rect 86310 2456 86316 2508
rect 86368 2496 86374 2508
rect 89530 2496 89536 2508
rect 86368 2468 89536 2496
rect 86368 2456 86374 2468
rect 89530 2456 89536 2468
rect 89588 2456 89594 2508
rect 91020 2468 110000 2496
rect 81544 2400 81664 2428
rect 76285 2363 76343 2369
rect 76285 2329 76297 2363
rect 76331 2360 76343 2363
rect 77021 2363 77079 2369
rect 77021 2360 77033 2363
rect 76331 2332 77033 2360
rect 76331 2329 76343 2332
rect 76285 2323 76343 2329
rect 77021 2329 77033 2332
rect 77067 2360 77079 2363
rect 81526 2360 81532 2372
rect 77067 2332 81532 2360
rect 77067 2329 77079 2332
rect 77021 2323 77079 2329
rect 81526 2320 81532 2332
rect 81584 2320 81590 2372
rect 81636 2360 81664 2400
rect 81986 2388 81992 2440
rect 82044 2428 82050 2440
rect 82357 2431 82415 2437
rect 82357 2428 82369 2431
rect 82044 2400 82369 2428
rect 82044 2388 82050 2400
rect 82357 2397 82369 2400
rect 82403 2397 82415 2431
rect 82357 2391 82415 2397
rect 83090 2388 83096 2440
rect 83148 2428 83154 2440
rect 83645 2431 83703 2437
rect 83645 2428 83657 2431
rect 83148 2400 83657 2428
rect 83148 2388 83154 2400
rect 83645 2397 83657 2400
rect 83691 2397 83703 2431
rect 84562 2428 84568 2440
rect 84523 2400 84568 2428
rect 83645 2391 83703 2397
rect 84562 2388 84568 2400
rect 84620 2388 84626 2440
rect 85298 2428 85304 2440
rect 85259 2400 85304 2428
rect 85298 2388 85304 2400
rect 85356 2388 85362 2440
rect 85666 2388 85672 2440
rect 85724 2428 85730 2440
rect 86405 2431 86463 2437
rect 86405 2428 86417 2431
rect 85724 2400 86417 2428
rect 85724 2388 85730 2400
rect 86405 2397 86417 2400
rect 86451 2397 86463 2431
rect 86405 2391 86463 2397
rect 87417 2431 87475 2437
rect 87417 2397 87429 2431
rect 87463 2428 87475 2431
rect 87598 2428 87604 2440
rect 87463 2400 87604 2428
rect 87463 2397 87475 2400
rect 87417 2391 87475 2397
rect 87598 2388 87604 2400
rect 87656 2388 87662 2440
rect 87690 2388 87696 2440
rect 87748 2428 87754 2440
rect 87748 2400 87793 2428
rect 87748 2388 87754 2400
rect 88978 2388 88984 2440
rect 89036 2428 89042 2440
rect 89036 2400 89081 2428
rect 89036 2388 89042 2400
rect 89162 2388 89168 2440
rect 89220 2428 89226 2440
rect 89809 2431 89867 2437
rect 89809 2428 89821 2431
rect 89220 2400 89821 2428
rect 89220 2388 89226 2400
rect 89809 2397 89821 2400
rect 89855 2397 89867 2431
rect 90450 2428 90456 2440
rect 90411 2400 90456 2428
rect 89809 2391 89867 2397
rect 90450 2388 90456 2400
rect 90508 2388 90514 2440
rect 81636 2332 82032 2360
rect 76561 2295 76619 2301
rect 76561 2292 76573 2295
rect 75656 2264 76573 2292
rect 75549 2255 75607 2261
rect 76561 2261 76573 2264
rect 76607 2261 76619 2295
rect 76561 2255 76619 2261
rect 76834 2252 76840 2304
rect 76892 2292 76898 2304
rect 76929 2295 76987 2301
rect 76929 2292 76941 2295
rect 76892 2264 76941 2292
rect 76892 2252 76898 2264
rect 76929 2261 76941 2264
rect 76975 2261 76987 2295
rect 76929 2255 76987 2261
rect 77110 2252 77116 2304
rect 77168 2292 77174 2304
rect 77386 2292 77392 2304
rect 77168 2264 77392 2292
rect 77168 2252 77174 2264
rect 77386 2252 77392 2264
rect 77444 2252 77450 2304
rect 77754 2292 77760 2304
rect 77715 2264 77760 2292
rect 77754 2252 77760 2264
rect 77812 2252 77818 2304
rect 78582 2252 78588 2304
rect 78640 2292 78646 2304
rect 78677 2295 78735 2301
rect 78677 2292 78689 2295
rect 78640 2264 78689 2292
rect 78640 2252 78646 2264
rect 78677 2261 78689 2264
rect 78723 2261 78735 2295
rect 78677 2255 78735 2261
rect 79226 2252 79232 2304
rect 79284 2292 79290 2304
rect 79321 2295 79379 2301
rect 79321 2292 79333 2295
rect 79284 2264 79333 2292
rect 79284 2252 79290 2264
rect 79321 2261 79333 2264
rect 79367 2261 79379 2295
rect 82004 2292 82032 2332
rect 82078 2320 82084 2372
rect 82136 2360 82142 2372
rect 91020 2360 91048 2468
rect 91462 2388 91468 2440
rect 91520 2428 91526 2440
rect 91741 2431 91799 2437
rect 91741 2428 91753 2431
rect 91520 2400 91753 2428
rect 91520 2388 91526 2400
rect 91741 2397 91753 2400
rect 91787 2397 91799 2431
rect 91741 2391 91799 2397
rect 92106 2388 92112 2440
rect 92164 2428 92170 2440
rect 92385 2431 92443 2437
rect 92385 2428 92397 2431
rect 92164 2400 92397 2428
rect 92164 2388 92170 2400
rect 92385 2397 92397 2400
rect 92431 2397 92443 2431
rect 92385 2391 92443 2397
rect 92750 2388 92756 2440
rect 92808 2428 92814 2440
rect 92845 2431 92903 2437
rect 92845 2428 92857 2431
rect 92808 2400 92857 2428
rect 92808 2388 92814 2400
rect 92845 2397 92857 2400
rect 92891 2397 92903 2431
rect 94314 2428 94320 2440
rect 94275 2400 94320 2428
rect 92845 2391 92903 2397
rect 94314 2388 94320 2400
rect 94372 2388 94378 2440
rect 95973 2431 96031 2437
rect 95973 2428 95985 2431
rect 94424 2400 95985 2428
rect 82136 2332 91048 2360
rect 82136 2320 82142 2332
rect 92290 2320 92296 2372
rect 92348 2360 92354 2372
rect 94424 2360 94452 2400
rect 95973 2397 95985 2400
rect 96019 2397 96031 2431
rect 95973 2391 96031 2397
rect 99650 2388 99656 2440
rect 99708 2428 99714 2440
rect 99745 2431 99803 2437
rect 99745 2428 99757 2431
rect 99708 2400 99757 2428
rect 99708 2388 99714 2400
rect 99745 2397 99757 2400
rect 99791 2397 99803 2431
rect 99745 2391 99803 2397
rect 100478 2388 100484 2440
rect 100536 2428 100542 2440
rect 100573 2431 100631 2437
rect 100573 2428 100585 2431
rect 100536 2400 100585 2428
rect 100536 2388 100542 2400
rect 100573 2397 100585 2400
rect 100619 2397 100631 2431
rect 100573 2391 100631 2397
rect 100662 2388 100668 2440
rect 100720 2428 100726 2440
rect 104526 2428 104532 2440
rect 100720 2400 104532 2428
rect 100720 2388 100726 2400
rect 104526 2388 104532 2400
rect 104584 2388 104590 2440
rect 104621 2431 104679 2437
rect 104621 2397 104633 2431
rect 104667 2428 104679 2431
rect 104894 2428 104900 2440
rect 104667 2400 104900 2428
rect 104667 2397 104679 2400
rect 104621 2391 104679 2397
rect 104894 2388 104900 2400
rect 104952 2388 104958 2440
rect 105998 2428 106004 2440
rect 105959 2400 106004 2428
rect 105998 2388 106004 2400
rect 106056 2388 106062 2440
rect 107013 2431 107071 2437
rect 107013 2397 107025 2431
rect 107059 2428 107071 2431
rect 107470 2428 107476 2440
rect 107059 2400 107476 2428
rect 107059 2397 107071 2400
rect 107013 2391 107071 2397
rect 107470 2388 107476 2400
rect 107528 2388 107534 2440
rect 107657 2431 107715 2437
rect 107657 2397 107669 2431
rect 107703 2397 107715 2431
rect 107657 2391 107715 2397
rect 92348 2332 94452 2360
rect 92348 2320 92354 2332
rect 94682 2320 94688 2372
rect 94740 2360 94746 2372
rect 94869 2363 94927 2369
rect 94869 2360 94881 2363
rect 94740 2332 94881 2360
rect 94740 2320 94746 2332
rect 94869 2329 94881 2332
rect 94915 2329 94927 2363
rect 94869 2323 94927 2329
rect 96614 2320 96620 2372
rect 96672 2360 96678 2372
rect 96985 2363 97043 2369
rect 96985 2360 96997 2363
rect 96672 2332 96997 2360
rect 96672 2320 96678 2332
rect 96985 2329 96997 2332
rect 97031 2329 97043 2363
rect 96985 2323 97043 2329
rect 97902 2320 97908 2372
rect 97960 2360 97966 2372
rect 98089 2363 98147 2369
rect 98089 2360 98101 2363
rect 97960 2332 98101 2360
rect 97960 2320 97966 2332
rect 98089 2329 98101 2332
rect 98135 2329 98147 2363
rect 98089 2323 98147 2329
rect 99190 2320 99196 2372
rect 99248 2360 99254 2372
rect 99561 2363 99619 2369
rect 99561 2360 99573 2363
rect 99248 2332 99573 2360
rect 99248 2320 99254 2332
rect 99561 2329 99573 2332
rect 99607 2329 99619 2363
rect 99561 2323 99619 2329
rect 101122 2320 101128 2372
rect 101180 2360 101186 2372
rect 102137 2363 102195 2369
rect 102137 2360 102149 2363
rect 101180 2332 102149 2360
rect 101180 2320 101186 2332
rect 102137 2329 102149 2332
rect 102183 2329 102195 2363
rect 102137 2323 102195 2329
rect 103054 2320 103060 2372
rect 103112 2360 103118 2372
rect 103241 2363 103299 2369
rect 103241 2360 103253 2363
rect 103112 2332 103253 2360
rect 103112 2320 103118 2332
rect 103241 2329 103253 2332
rect 103287 2329 103299 2363
rect 103241 2323 103299 2329
rect 104986 2320 104992 2372
rect 105044 2360 105050 2372
rect 105173 2363 105231 2369
rect 105173 2360 105185 2363
rect 105044 2332 105185 2360
rect 105044 2320 105050 2332
rect 105173 2329 105185 2332
rect 105219 2329 105231 2363
rect 107672 2360 107700 2391
rect 108114 2388 108120 2440
rect 108172 2388 108178 2440
rect 108298 2388 108304 2440
rect 108356 2428 108362 2440
rect 108356 2400 108401 2428
rect 108356 2388 108362 2400
rect 105173 2323 105231 2329
rect 106844 2332 107700 2360
rect 83829 2295 83887 2301
rect 83829 2292 83841 2295
rect 82004 2264 83841 2292
rect 79321 2255 79379 2261
rect 83829 2261 83841 2264
rect 83875 2261 83887 2295
rect 83829 2255 83887 2261
rect 84010 2252 84016 2304
rect 84068 2292 84074 2304
rect 84381 2295 84439 2301
rect 84381 2292 84393 2295
rect 84068 2264 84393 2292
rect 84068 2252 84074 2264
rect 84381 2261 84393 2264
rect 84427 2261 84439 2295
rect 84381 2255 84439 2261
rect 85022 2252 85028 2304
rect 85080 2292 85086 2304
rect 85117 2295 85175 2301
rect 85117 2292 85129 2295
rect 85080 2264 85129 2292
rect 85080 2252 85086 2264
rect 85117 2261 85129 2264
rect 85163 2261 85175 2295
rect 85117 2255 85175 2261
rect 85482 2252 85488 2304
rect 85540 2292 85546 2304
rect 86221 2295 86279 2301
rect 86221 2292 86233 2295
rect 85540 2264 86233 2292
rect 85540 2252 85546 2264
rect 86221 2261 86233 2264
rect 86267 2261 86279 2295
rect 86221 2255 86279 2261
rect 88242 2252 88248 2304
rect 88300 2292 88306 2304
rect 88797 2295 88855 2301
rect 88797 2292 88809 2295
rect 88300 2264 88809 2292
rect 88300 2252 88306 2264
rect 88797 2261 88809 2264
rect 88843 2261 88855 2295
rect 88797 2255 88855 2261
rect 89162 2252 89168 2304
rect 89220 2292 89226 2304
rect 89625 2295 89683 2301
rect 89625 2292 89637 2295
rect 89220 2264 89637 2292
rect 89220 2252 89226 2264
rect 89625 2261 89637 2264
rect 89671 2261 89683 2295
rect 89625 2255 89683 2261
rect 90174 2252 90180 2304
rect 90232 2292 90238 2304
rect 90269 2295 90327 2301
rect 90269 2292 90281 2295
rect 90232 2264 90281 2292
rect 90232 2252 90238 2264
rect 90269 2261 90281 2264
rect 90315 2261 90327 2295
rect 91554 2292 91560 2304
rect 91515 2264 91560 2292
rect 90269 2255 90327 2261
rect 91554 2252 91560 2264
rect 91612 2252 91618 2304
rect 92198 2292 92204 2304
rect 92159 2264 92204 2292
rect 92198 2252 92204 2264
rect 92256 2252 92262 2304
rect 93026 2292 93032 2304
rect 92987 2264 93032 2292
rect 93026 2252 93032 2264
rect 93084 2252 93090 2304
rect 94038 2252 94044 2304
rect 94096 2292 94102 2304
rect 94133 2295 94191 2301
rect 94133 2292 94145 2295
rect 94096 2264 94145 2292
rect 94096 2252 94102 2264
rect 94133 2261 94145 2264
rect 94179 2261 94191 2295
rect 94958 2292 94964 2304
rect 94919 2264 94964 2292
rect 94133 2255 94191 2261
rect 94958 2252 94964 2264
rect 95016 2252 95022 2304
rect 95789 2295 95847 2301
rect 95789 2261 95801 2295
rect 95835 2292 95847 2295
rect 95970 2292 95976 2304
rect 95835 2264 95976 2292
rect 95835 2261 95847 2264
rect 95789 2255 95847 2261
rect 95970 2252 95976 2264
rect 96028 2252 96034 2304
rect 97074 2292 97080 2304
rect 97035 2264 97080 2292
rect 97074 2252 97080 2264
rect 97132 2252 97138 2304
rect 98178 2292 98184 2304
rect 98139 2264 98184 2292
rect 98178 2252 98184 2264
rect 98236 2252 98242 2304
rect 104342 2252 104348 2304
rect 104400 2292 104406 2304
rect 104437 2295 104495 2301
rect 104437 2292 104449 2295
rect 104400 2264 104449 2292
rect 104400 2252 104406 2264
rect 104437 2261 104449 2264
rect 104483 2261 104495 2295
rect 105262 2292 105268 2304
rect 105223 2264 105268 2292
rect 104437 2255 104495 2261
rect 105262 2252 105268 2264
rect 105320 2252 105326 2304
rect 105630 2252 105636 2304
rect 105688 2292 105694 2304
rect 106844 2301 106872 2332
rect 105817 2295 105875 2301
rect 105817 2292 105829 2295
rect 105688 2264 105829 2292
rect 105688 2252 105694 2264
rect 105817 2261 105829 2264
rect 105863 2261 105875 2295
rect 105817 2255 105875 2261
rect 106829 2295 106887 2301
rect 106829 2261 106841 2295
rect 106875 2261 106887 2295
rect 106829 2255 106887 2261
rect 106918 2252 106924 2304
rect 106976 2292 106982 2304
rect 108132 2301 108160 2388
rect 108850 2320 108856 2372
rect 108908 2360 108914 2372
rect 109865 2363 109923 2369
rect 109865 2360 109877 2363
rect 108908 2332 109877 2360
rect 108908 2320 108914 2332
rect 109865 2329 109877 2332
rect 109911 2329 109923 2363
rect 109972 2360 110000 2468
rect 110046 2456 110052 2508
rect 110104 2496 110110 2508
rect 117869 2499 117927 2505
rect 117869 2496 117881 2499
rect 110104 2468 117881 2496
rect 110104 2456 110110 2468
rect 117869 2465 117881 2468
rect 117915 2465 117927 2499
rect 117869 2459 117927 2465
rect 110782 2388 110788 2440
rect 110840 2428 110846 2440
rect 110877 2431 110935 2437
rect 110877 2428 110889 2431
rect 110840 2400 110889 2428
rect 110840 2388 110846 2400
rect 110877 2397 110889 2400
rect 110923 2397 110935 2431
rect 110877 2391 110935 2397
rect 112070 2388 112076 2440
rect 112128 2428 112134 2440
rect 112165 2431 112223 2437
rect 112165 2428 112177 2431
rect 112128 2400 112177 2428
rect 112128 2388 112134 2400
rect 112165 2397 112177 2400
rect 112211 2397 112223 2431
rect 112438 2428 112444 2440
rect 112399 2400 112444 2428
rect 112165 2391 112223 2397
rect 112438 2388 112444 2400
rect 112496 2388 112502 2440
rect 113634 2428 113640 2440
rect 113595 2400 113640 2428
rect 113634 2388 113640 2400
rect 113692 2388 113698 2440
rect 114002 2388 114008 2440
rect 114060 2428 114066 2440
rect 114741 2431 114799 2437
rect 114741 2428 114753 2431
rect 114060 2400 114753 2428
rect 114060 2388 114066 2400
rect 114741 2397 114753 2400
rect 114787 2397 114799 2431
rect 114741 2391 114799 2397
rect 115290 2388 115296 2440
rect 115348 2428 115354 2440
rect 115385 2431 115443 2437
rect 115385 2428 115397 2431
rect 115348 2400 115397 2428
rect 115348 2388 115354 2400
rect 115385 2397 115397 2400
rect 115431 2397 115443 2431
rect 118142 2428 118148 2440
rect 115385 2391 115443 2397
rect 115676 2400 118148 2428
rect 115676 2360 115704 2400
rect 118142 2388 118148 2400
rect 118200 2388 118206 2440
rect 116394 2360 116400 2372
rect 109972 2332 115704 2360
rect 116355 2332 116400 2360
rect 109865 2323 109923 2329
rect 116394 2320 116400 2332
rect 116452 2320 116458 2372
rect 116578 2320 116584 2372
rect 116636 2360 116642 2372
rect 117593 2363 117651 2369
rect 117593 2360 117605 2363
rect 116636 2332 117605 2360
rect 116636 2320 116642 2332
rect 117593 2329 117605 2332
rect 117639 2329 117651 2363
rect 117593 2323 117651 2329
rect 107473 2295 107531 2301
rect 107473 2292 107485 2295
rect 106976 2264 107485 2292
rect 106976 2252 106982 2264
rect 107473 2261 107485 2264
rect 107519 2261 107531 2295
rect 107473 2255 107531 2261
rect 108117 2295 108175 2301
rect 108117 2261 108129 2295
rect 108163 2261 108175 2295
rect 109954 2292 109960 2304
rect 109915 2264 109960 2292
rect 108117 2255 108175 2261
rect 109954 2252 109960 2264
rect 110012 2252 110018 2304
rect 113358 2252 113364 2304
rect 113416 2292 113422 2304
rect 113453 2295 113511 2301
rect 113453 2292 113465 2295
rect 113416 2264 113465 2292
rect 113416 2252 113422 2264
rect 113453 2261 113465 2264
rect 113499 2261 113511 2295
rect 115566 2292 115572 2304
rect 115527 2264 115572 2292
rect 113453 2255 113511 2261
rect 115566 2252 115572 2264
rect 115624 2252 115630 2304
rect 116486 2292 116492 2304
rect 116447 2264 116492 2292
rect 116486 2252 116492 2264
rect 116544 2252 116550 2304
rect 1104 2202 118864 2224
rect 1104 2150 30398 2202
rect 30450 2150 30462 2202
rect 30514 2150 30526 2202
rect 30578 2150 30590 2202
rect 30642 2150 30654 2202
rect 30706 2150 59846 2202
rect 59898 2150 59910 2202
rect 59962 2150 59974 2202
rect 60026 2150 60038 2202
rect 60090 2150 60102 2202
rect 60154 2150 89294 2202
rect 89346 2150 89358 2202
rect 89410 2150 89422 2202
rect 89474 2150 89486 2202
rect 89538 2150 89550 2202
rect 89602 2150 118864 2202
rect 1104 2128 118864 2150
rect 10134 2048 10140 2100
rect 10192 2088 10198 2100
rect 60642 2088 60648 2100
rect 10192 2060 60648 2088
rect 10192 2048 10198 2060
rect 60642 2048 60648 2060
rect 60700 2048 60706 2100
rect 60734 2048 60740 2100
rect 60792 2088 60798 2100
rect 66070 2088 66076 2100
rect 60792 2060 66076 2088
rect 60792 2048 60798 2060
rect 66070 2048 66076 2060
rect 66128 2048 66134 2100
rect 66806 2048 66812 2100
rect 66864 2088 66870 2100
rect 66864 2060 67128 2088
rect 66864 2048 66870 2060
rect 1670 1980 1676 2032
rect 1728 2020 1734 2032
rect 28258 2020 28264 2032
rect 1728 1992 28264 2020
rect 1728 1980 1734 1992
rect 28258 1980 28264 1992
rect 28316 1980 28322 2032
rect 28442 1980 28448 2032
rect 28500 2020 28506 2032
rect 29822 2020 29828 2032
rect 28500 1992 29828 2020
rect 28500 1980 28506 1992
rect 29822 1980 29828 1992
rect 29880 1980 29886 2032
rect 30742 1980 30748 2032
rect 30800 2020 30806 2032
rect 37734 2020 37740 2032
rect 30800 1992 37740 2020
rect 30800 1980 30806 1992
rect 37734 1980 37740 1992
rect 37792 1980 37798 2032
rect 38654 1980 38660 2032
rect 38712 2020 38718 2032
rect 60918 2020 60924 2032
rect 38712 1992 60924 2020
rect 38712 1980 38718 1992
rect 60918 1980 60924 1992
rect 60976 1980 60982 2032
rect 61010 1980 61016 2032
rect 61068 2020 61074 2032
rect 63494 2020 63500 2032
rect 61068 1992 63500 2020
rect 61068 1980 61074 1992
rect 63494 1980 63500 1992
rect 63552 1980 63558 2032
rect 67100 2020 67128 2060
rect 67174 2048 67180 2100
rect 67232 2088 67238 2100
rect 73522 2088 73528 2100
rect 67232 2060 73528 2088
rect 67232 2048 67238 2060
rect 73522 2048 73528 2060
rect 73580 2048 73586 2100
rect 73614 2048 73620 2100
rect 73672 2088 73678 2100
rect 118050 2088 118056 2100
rect 73672 2060 118056 2088
rect 73672 2048 73678 2060
rect 118050 2048 118056 2060
rect 118108 2048 118114 2100
rect 116486 2020 116492 2032
rect 67100 1992 116492 2020
rect 116486 1980 116492 1992
rect 116544 1980 116550 2032
rect 12526 1912 12532 1964
rect 12584 1952 12590 1964
rect 40494 1952 40500 1964
rect 12584 1924 40500 1952
rect 12584 1912 12590 1924
rect 40494 1912 40500 1924
rect 40552 1912 40558 1964
rect 40862 1912 40868 1964
rect 40920 1952 40926 1964
rect 40920 1924 45554 1952
rect 40920 1912 40926 1924
rect 7374 1844 7380 1896
rect 7432 1884 7438 1896
rect 31386 1884 31392 1896
rect 7432 1856 31392 1884
rect 7432 1844 7438 1856
rect 31386 1844 31392 1856
rect 31444 1844 31450 1896
rect 31570 1844 31576 1896
rect 31628 1884 31634 1896
rect 38470 1884 38476 1896
rect 31628 1856 38476 1884
rect 31628 1844 31634 1856
rect 38470 1844 38476 1856
rect 38528 1844 38534 1896
rect 45526 1884 45554 1924
rect 46658 1912 46664 1964
rect 46716 1952 46722 1964
rect 55214 1952 55220 1964
rect 46716 1924 55220 1952
rect 46716 1912 46722 1924
rect 55214 1912 55220 1924
rect 55272 1912 55278 1964
rect 55306 1912 55312 1964
rect 55364 1952 55370 1964
rect 60734 1952 60740 1964
rect 55364 1924 60740 1952
rect 55364 1912 55370 1924
rect 60734 1912 60740 1924
rect 60792 1912 60798 1964
rect 60826 1912 60832 1964
rect 60884 1952 60890 1964
rect 73890 1952 73896 1964
rect 60884 1924 73896 1952
rect 60884 1912 60890 1924
rect 73890 1912 73896 1924
rect 73948 1912 73954 1964
rect 73982 1912 73988 1964
rect 74040 1952 74046 1964
rect 105262 1952 105268 1964
rect 74040 1924 105268 1952
rect 74040 1912 74046 1924
rect 105262 1912 105268 1924
rect 105320 1912 105326 1964
rect 70946 1884 70952 1896
rect 45526 1856 70952 1884
rect 70946 1844 70952 1856
rect 71004 1844 71010 1896
rect 71038 1844 71044 1896
rect 71096 1884 71102 1896
rect 75362 1884 75368 1896
rect 71096 1856 75368 1884
rect 71096 1844 71102 1856
rect 75362 1844 75368 1856
rect 75420 1844 75426 1896
rect 75546 1844 75552 1896
rect 75604 1884 75610 1896
rect 77202 1884 77208 1896
rect 75604 1856 77208 1884
rect 75604 1844 75610 1856
rect 77202 1844 77208 1856
rect 77260 1844 77266 1896
rect 77386 1844 77392 1896
rect 77444 1884 77450 1896
rect 109770 1884 109776 1896
rect 77444 1856 109776 1884
rect 77444 1844 77450 1856
rect 109770 1844 109776 1856
rect 109828 1844 109834 1896
rect 15746 1776 15752 1828
rect 15804 1816 15810 1828
rect 42702 1816 42708 1828
rect 15804 1788 42708 1816
rect 15804 1776 15810 1788
rect 42702 1776 42708 1788
rect 42760 1776 42766 1828
rect 45922 1776 45928 1828
rect 45980 1816 45986 1828
rect 45980 1788 49832 1816
rect 45980 1776 45986 1788
rect 17494 1708 17500 1760
rect 17552 1748 17558 1760
rect 27706 1748 27712 1760
rect 17552 1720 27712 1748
rect 17552 1708 17558 1720
rect 27706 1708 27712 1720
rect 27764 1708 27770 1760
rect 29730 1708 29736 1760
rect 29788 1748 29794 1760
rect 49694 1748 49700 1760
rect 29788 1720 49700 1748
rect 29788 1708 29794 1720
rect 49694 1708 49700 1720
rect 49752 1708 49758 1760
rect 49804 1748 49832 1788
rect 51534 1776 51540 1828
rect 51592 1816 51598 1828
rect 58158 1816 58164 1828
rect 51592 1788 58164 1816
rect 51592 1776 51598 1788
rect 58158 1776 58164 1788
rect 58216 1776 58222 1828
rect 58250 1776 58256 1828
rect 58308 1816 58314 1828
rect 89530 1816 89536 1828
rect 58308 1788 89536 1816
rect 58308 1776 58314 1788
rect 89530 1776 89536 1788
rect 89588 1776 89594 1828
rect 89622 1776 89628 1828
rect 89680 1816 89686 1828
rect 89680 1788 94544 1816
rect 89680 1776 89686 1788
rect 51626 1748 51632 1760
rect 49804 1720 51632 1748
rect 51626 1708 51632 1720
rect 51684 1708 51690 1760
rect 51810 1708 51816 1760
rect 51868 1748 51874 1760
rect 51868 1720 75224 1748
rect 51868 1708 51874 1720
rect 3510 1640 3516 1692
rect 3568 1680 3574 1692
rect 55950 1680 55956 1692
rect 3568 1652 55956 1680
rect 3568 1640 3574 1652
rect 55950 1640 55956 1652
rect 56008 1640 56014 1692
rect 56410 1640 56416 1692
rect 56468 1680 56474 1692
rect 58066 1680 58072 1692
rect 56468 1652 58072 1680
rect 56468 1640 56474 1652
rect 58066 1640 58072 1652
rect 58124 1640 58130 1692
rect 66898 1640 66904 1692
rect 66956 1680 66962 1692
rect 71314 1680 71320 1692
rect 66956 1652 71320 1680
rect 66956 1640 66962 1652
rect 71314 1640 71320 1652
rect 71372 1640 71378 1692
rect 71866 1640 71872 1692
rect 71924 1680 71930 1692
rect 73982 1680 73988 1692
rect 71924 1652 73988 1680
rect 71924 1640 71930 1652
rect 73982 1640 73988 1652
rect 74040 1640 74046 1692
rect 74074 1640 74080 1692
rect 74132 1680 74138 1692
rect 75086 1680 75092 1692
rect 74132 1652 75092 1680
rect 74132 1640 74138 1652
rect 75086 1640 75092 1652
rect 75144 1640 75150 1692
rect 75196 1680 75224 1720
rect 76834 1708 76840 1760
rect 76892 1748 76898 1760
rect 91554 1748 91560 1760
rect 76892 1720 91560 1748
rect 76892 1708 76898 1720
rect 91554 1708 91560 1720
rect 91612 1708 91618 1760
rect 94516 1748 94544 1788
rect 94774 1776 94780 1828
rect 94832 1816 94838 1828
rect 94832 1788 100800 1816
rect 94832 1776 94838 1788
rect 100662 1748 100668 1760
rect 94516 1720 100668 1748
rect 100662 1708 100668 1720
rect 100720 1708 100726 1760
rect 100772 1748 100800 1788
rect 100846 1776 100852 1828
rect 100904 1816 100910 1828
rect 105998 1816 106004 1828
rect 100904 1788 106004 1816
rect 100904 1776 100910 1788
rect 105998 1776 106004 1788
rect 106056 1776 106062 1828
rect 112438 1748 112444 1760
rect 100772 1720 112444 1748
rect 112438 1708 112444 1720
rect 112496 1708 112502 1760
rect 77754 1680 77760 1692
rect 75196 1652 77760 1680
rect 77754 1640 77760 1652
rect 77812 1640 77818 1692
rect 77846 1640 77852 1692
rect 77904 1680 77910 1692
rect 98178 1680 98184 1692
rect 77904 1652 98184 1680
rect 77904 1640 77910 1652
rect 98178 1640 98184 1652
rect 98236 1640 98242 1692
rect 7190 1572 7196 1624
rect 7248 1612 7254 1624
rect 45554 1612 45560 1624
rect 7248 1584 45560 1612
rect 7248 1572 7254 1584
rect 45554 1572 45560 1584
rect 45612 1572 45618 1624
rect 45646 1572 45652 1624
rect 45704 1612 45710 1624
rect 51994 1612 52000 1624
rect 45704 1584 52000 1612
rect 45704 1572 45710 1584
rect 51994 1572 52000 1584
rect 52052 1572 52058 1624
rect 53098 1572 53104 1624
rect 53156 1612 53162 1624
rect 109954 1612 109960 1624
rect 53156 1584 109960 1612
rect 53156 1572 53162 1584
rect 109954 1572 109960 1584
rect 110012 1572 110018 1624
rect 12342 1504 12348 1556
rect 12400 1544 12406 1556
rect 12400 1516 89576 1544
rect 12400 1504 12406 1516
rect 18230 1436 18236 1488
rect 18288 1476 18294 1488
rect 30742 1476 30748 1488
rect 18288 1448 30748 1476
rect 18288 1436 18294 1448
rect 30742 1436 30748 1448
rect 30800 1436 30806 1488
rect 31662 1436 31668 1488
rect 31720 1476 31726 1488
rect 89346 1476 89352 1488
rect 31720 1448 89352 1476
rect 31720 1436 31726 1448
rect 89346 1436 89352 1448
rect 89404 1436 89410 1488
rect 89548 1476 89576 1516
rect 89622 1504 89628 1556
rect 89680 1544 89686 1556
rect 89714 1544 89720 1556
rect 89680 1516 89720 1544
rect 89680 1504 89686 1516
rect 89714 1504 89720 1516
rect 89772 1504 89778 1556
rect 89806 1504 89812 1556
rect 89864 1544 89870 1556
rect 94314 1544 94320 1556
rect 89864 1516 94320 1544
rect 89864 1504 89870 1516
rect 94314 1504 94320 1516
rect 94372 1504 94378 1556
rect 97810 1504 97816 1556
rect 97868 1544 97874 1556
rect 100846 1544 100852 1556
rect 97868 1516 100852 1544
rect 97868 1504 97874 1516
rect 100846 1504 100852 1516
rect 100904 1504 100910 1556
rect 94958 1476 94964 1488
rect 89548 1448 94964 1476
rect 94958 1436 94964 1448
rect 95016 1436 95022 1488
rect 7006 1368 7012 1420
rect 7064 1408 7070 1420
rect 80054 1408 80060 1420
rect 7064 1380 80060 1408
rect 7064 1368 7070 1380
rect 80054 1368 80060 1380
rect 80112 1368 80118 1420
rect 80146 1368 80152 1420
rect 80204 1408 80210 1420
rect 86494 1408 86500 1420
rect 80204 1380 86500 1408
rect 80204 1368 80210 1380
rect 86494 1368 86500 1380
rect 86552 1368 86558 1420
rect 86586 1368 86592 1420
rect 86644 1408 86650 1420
rect 89438 1408 89444 1420
rect 86644 1380 89444 1408
rect 86644 1368 86650 1380
rect 89438 1368 89444 1380
rect 89496 1368 89502 1420
rect 89530 1368 89536 1420
rect 89588 1408 89594 1420
rect 97074 1408 97080 1420
rect 89588 1380 97080 1408
rect 89588 1368 89594 1380
rect 97074 1368 97080 1380
rect 97132 1368 97138 1420
rect 107562 1368 107568 1420
rect 107620 1408 107626 1420
rect 108298 1408 108304 1420
rect 107620 1380 108304 1408
rect 107620 1368 107626 1380
rect 108298 1368 108304 1380
rect 108356 1368 108362 1420
rect 28902 1300 28908 1352
rect 28960 1340 28966 1352
rect 93026 1340 93032 1352
rect 28960 1312 93032 1340
rect 28960 1300 28966 1312
rect 93026 1300 93032 1312
rect 93084 1300 93090 1352
rect 22462 1232 22468 1284
rect 22520 1272 22526 1284
rect 31662 1272 31668 1284
rect 22520 1244 31668 1272
rect 22520 1232 22526 1244
rect 31662 1232 31668 1244
rect 31720 1232 31726 1284
rect 41782 1232 41788 1284
rect 41840 1272 41846 1284
rect 90450 1272 90456 1284
rect 41840 1244 90456 1272
rect 41840 1232 41846 1244
rect 90450 1232 90456 1244
rect 90508 1232 90514 1284
rect 47946 1164 47952 1216
rect 48004 1204 48010 1216
rect 81342 1204 81348 1216
rect 48004 1176 81348 1204
rect 48004 1164 48010 1176
rect 81342 1164 81348 1176
rect 81400 1164 81406 1216
rect 86494 1164 86500 1216
rect 86552 1204 86558 1216
rect 89530 1204 89536 1216
rect 86552 1176 89536 1204
rect 86552 1164 86558 1176
rect 89530 1164 89536 1176
rect 89588 1164 89594 1216
rect 57146 1096 57152 1148
rect 57204 1136 57210 1148
rect 87690 1136 87696 1148
rect 57204 1108 87696 1136
rect 57204 1096 57210 1108
rect 87690 1096 87696 1108
rect 87748 1096 87754 1148
<< via1 >>
rect 50804 28092 50856 28144
rect 53104 28092 53156 28144
rect 40868 28024 40920 28076
rect 46756 28024 46808 28076
rect 50712 28024 50764 28076
rect 57612 28024 57664 28076
rect 69296 28024 69348 28076
rect 75276 28024 75328 28076
rect 26700 27956 26752 28008
rect 39580 27956 39632 28008
rect 39672 27956 39724 28008
rect 40408 27956 40460 28008
rect 49148 27956 49200 28008
rect 49700 27956 49752 28008
rect 50252 27956 50304 28008
rect 53472 27956 53524 28008
rect 59084 27956 59136 28008
rect 62948 27956 63000 28008
rect 70308 27956 70360 28008
rect 75000 27956 75052 28008
rect 9864 27820 9916 27872
rect 17132 27820 17184 27872
rect 19800 27820 19852 27872
rect 27068 27820 27120 27872
rect 31760 27820 31812 27872
rect 40868 27888 40920 27940
rect 40960 27888 41012 27940
rect 41420 27888 41472 27940
rect 46480 27888 46532 27940
rect 59728 27888 59780 27940
rect 61476 27888 61528 27940
rect 68744 27888 68796 27940
rect 72884 27888 72936 27940
rect 76196 27888 76248 27940
rect 32680 27820 32732 27872
rect 50804 27820 50856 27872
rect 50896 27820 50948 27872
rect 54668 27820 54720 27872
rect 59360 27820 59412 27872
rect 62120 27820 62172 27872
rect 68008 27820 68060 27872
rect 68928 27820 68980 27872
rect 74448 27820 74500 27872
rect 75920 27820 75972 27872
rect 78588 27820 78640 27872
rect 79600 27820 79652 27872
rect 79784 27820 79836 27872
rect 80428 27820 80480 27872
rect 84844 27820 84896 27872
rect 93676 27820 93728 27872
rect 15674 27718 15726 27770
rect 15738 27718 15790 27770
rect 15802 27718 15854 27770
rect 15866 27718 15918 27770
rect 15930 27718 15982 27770
rect 45122 27718 45174 27770
rect 45186 27718 45238 27770
rect 45250 27718 45302 27770
rect 45314 27718 45366 27770
rect 45378 27718 45430 27770
rect 74570 27718 74622 27770
rect 74634 27718 74686 27770
rect 74698 27718 74750 27770
rect 74762 27718 74814 27770
rect 74826 27718 74878 27770
rect 104018 27718 104070 27770
rect 104082 27718 104134 27770
rect 104146 27718 104198 27770
rect 104210 27718 104262 27770
rect 104274 27718 104326 27770
rect 17132 27616 17184 27668
rect 84844 27616 84896 27668
rect 89720 27616 89772 27668
rect 101680 27659 101732 27668
rect 9588 27548 9640 27600
rect 9864 27548 9916 27600
rect 17040 27548 17092 27600
rect 18696 27548 18748 27600
rect 19340 27548 19392 27600
rect 22652 27591 22704 27600
rect 2412 27523 2464 27532
rect 2412 27489 2421 27523
rect 2421 27489 2455 27523
rect 2455 27489 2464 27523
rect 2412 27480 2464 27489
rect 4988 27523 5040 27532
rect 4988 27489 4997 27523
rect 4997 27489 5031 27523
rect 5031 27489 5040 27523
rect 4988 27480 5040 27489
rect 6368 27523 6420 27532
rect 6368 27489 6377 27523
rect 6377 27489 6411 27523
rect 6411 27489 6420 27523
rect 6368 27480 6420 27489
rect 22376 27480 22428 27532
rect 22652 27557 22661 27591
rect 22661 27557 22695 27591
rect 22695 27557 22704 27591
rect 22652 27548 22704 27557
rect 23388 27480 23440 27532
rect 2688 27455 2740 27464
rect 2688 27421 2697 27455
rect 2697 27421 2731 27455
rect 2731 27421 2740 27455
rect 2688 27412 2740 27421
rect 3608 27412 3660 27464
rect 6644 27455 6696 27464
rect 4436 27387 4488 27396
rect 4436 27353 4445 27387
rect 4445 27353 4479 27387
rect 4479 27353 4488 27387
rect 4436 27344 4488 27353
rect 1400 27319 1452 27328
rect 1400 27285 1409 27319
rect 1409 27285 1443 27319
rect 1443 27285 1452 27319
rect 1400 27276 1452 27285
rect 6644 27421 6653 27455
rect 6653 27421 6687 27455
rect 6687 27421 6696 27455
rect 6644 27412 6696 27421
rect 7104 27412 7156 27464
rect 11060 27412 11112 27464
rect 12440 27455 12492 27464
rect 12440 27421 12449 27455
rect 12449 27421 12483 27455
rect 12483 27421 12492 27455
rect 12440 27412 12492 27421
rect 13820 27412 13872 27464
rect 9404 27387 9456 27396
rect 9404 27353 9413 27387
rect 9413 27353 9447 27387
rect 9447 27353 9456 27387
rect 9404 27344 9456 27353
rect 10324 27387 10376 27396
rect 10324 27353 10333 27387
rect 10333 27353 10367 27387
rect 10367 27353 10376 27387
rect 10324 27344 10376 27353
rect 15200 27344 15252 27396
rect 16028 27412 16080 27464
rect 17224 27455 17276 27464
rect 17224 27421 17233 27455
rect 17233 27421 17267 27455
rect 17267 27421 17276 27455
rect 17224 27412 17276 27421
rect 18052 27412 18104 27464
rect 20168 27455 20220 27464
rect 16120 27344 16172 27396
rect 16212 27344 16264 27396
rect 19340 27344 19392 27396
rect 20168 27421 20177 27455
rect 20177 27421 20211 27455
rect 20211 27421 20220 27455
rect 20168 27412 20220 27421
rect 20352 27455 20404 27464
rect 20352 27421 20361 27455
rect 20361 27421 20395 27455
rect 20395 27421 20404 27455
rect 20352 27412 20404 27421
rect 20536 27412 20588 27464
rect 21088 27412 21140 27464
rect 21916 27344 21968 27396
rect 22100 27412 22152 27464
rect 27160 27548 27212 27600
rect 23572 27480 23624 27532
rect 23664 27412 23716 27464
rect 23848 27455 23900 27464
rect 23848 27421 23857 27455
rect 23857 27421 23891 27455
rect 23891 27421 23900 27455
rect 23848 27412 23900 27421
rect 25136 27412 25188 27464
rect 25320 27455 25372 27464
rect 25320 27421 25329 27455
rect 25329 27421 25363 27455
rect 25363 27421 25372 27455
rect 25320 27412 25372 27421
rect 26424 27412 26476 27464
rect 31392 27548 31444 27600
rect 11980 27276 12032 27328
rect 12532 27319 12584 27328
rect 12532 27285 12541 27319
rect 12541 27285 12575 27319
rect 12575 27285 12584 27319
rect 12532 27276 12584 27285
rect 17132 27276 17184 27328
rect 17316 27319 17368 27328
rect 17316 27285 17325 27319
rect 17325 27285 17359 27319
rect 17359 27285 17368 27319
rect 17316 27276 17368 27285
rect 20628 27276 20680 27328
rect 20812 27319 20864 27328
rect 20812 27285 20821 27319
rect 20821 27285 20855 27319
rect 20855 27285 20864 27319
rect 20812 27276 20864 27285
rect 22008 27319 22060 27328
rect 22008 27285 22017 27319
rect 22017 27285 22051 27319
rect 22051 27285 22060 27319
rect 22008 27276 22060 27285
rect 22284 27276 22336 27328
rect 23572 27276 23624 27328
rect 26884 27344 26936 27396
rect 27528 27344 27580 27396
rect 24400 27319 24452 27328
rect 24400 27285 24409 27319
rect 24409 27285 24443 27319
rect 24443 27285 24452 27319
rect 24400 27276 24452 27285
rect 26700 27276 26752 27328
rect 26976 27276 27028 27328
rect 30656 27480 30708 27532
rect 30748 27523 30800 27532
rect 30748 27489 30757 27523
rect 30757 27489 30791 27523
rect 30791 27489 30800 27523
rect 30748 27480 30800 27489
rect 31116 27480 31168 27532
rect 31760 27548 31812 27600
rect 28080 27455 28132 27464
rect 28080 27421 28089 27455
rect 28089 27421 28123 27455
rect 28123 27421 28132 27455
rect 28080 27412 28132 27421
rect 28908 27412 28960 27464
rect 30288 27344 30340 27396
rect 30840 27412 30892 27464
rect 30932 27412 30984 27464
rect 31852 27480 31904 27532
rect 33048 27548 33100 27600
rect 32036 27480 32088 27532
rect 33324 27523 33376 27532
rect 33324 27489 33333 27523
rect 33333 27489 33367 27523
rect 33367 27489 33376 27523
rect 33324 27480 33376 27489
rect 34704 27523 34756 27532
rect 31576 27344 31628 27396
rect 33600 27455 33652 27464
rect 32036 27344 32088 27396
rect 32128 27344 32180 27396
rect 33600 27421 33609 27455
rect 33609 27421 33643 27455
rect 33643 27421 33652 27455
rect 33600 27412 33652 27421
rect 34704 27489 34713 27523
rect 34713 27489 34747 27523
rect 34747 27489 34756 27523
rect 34704 27480 34756 27489
rect 34888 27548 34940 27600
rect 38200 27548 38252 27600
rect 39948 27548 40000 27600
rect 40592 27548 40644 27600
rect 40684 27548 40736 27600
rect 40408 27523 40460 27532
rect 40408 27489 40417 27523
rect 40417 27489 40451 27523
rect 40451 27489 40460 27523
rect 40408 27480 40460 27489
rect 41236 27480 41288 27532
rect 42800 27548 42852 27600
rect 43812 27480 43864 27532
rect 50528 27548 50580 27600
rect 53472 27591 53524 27600
rect 53472 27557 53481 27591
rect 53481 27557 53515 27591
rect 53515 27557 53524 27591
rect 53472 27548 53524 27557
rect 54116 27548 54168 27600
rect 59360 27548 59412 27600
rect 59452 27548 59504 27600
rect 61108 27548 61160 27600
rect 61200 27548 61252 27600
rect 34888 27412 34940 27464
rect 35072 27412 35124 27464
rect 32772 27387 32824 27396
rect 32772 27353 32781 27387
rect 32781 27353 32815 27387
rect 32815 27353 32824 27387
rect 32772 27344 32824 27353
rect 36268 27387 36320 27396
rect 36268 27353 36277 27387
rect 36277 27353 36311 27387
rect 36311 27353 36320 27387
rect 37372 27412 37424 27464
rect 39212 27412 39264 27464
rect 40500 27412 40552 27464
rect 40592 27412 40644 27464
rect 41880 27412 41932 27464
rect 43352 27455 43404 27464
rect 43352 27421 43361 27455
rect 43361 27421 43395 27455
rect 43395 27421 43404 27455
rect 43352 27412 43404 27421
rect 44088 27455 44140 27464
rect 44088 27421 44097 27455
rect 44097 27421 44131 27455
rect 44131 27421 44140 27455
rect 44088 27412 44140 27421
rect 44456 27412 44508 27464
rect 47216 27412 47268 27464
rect 48320 27412 48372 27464
rect 49148 27480 49200 27532
rect 54484 27523 54536 27532
rect 54484 27489 54493 27523
rect 54493 27489 54527 27523
rect 54527 27489 54536 27523
rect 54484 27480 54536 27489
rect 54668 27480 54720 27532
rect 60740 27480 60792 27532
rect 60924 27480 60976 27532
rect 36268 27344 36320 27353
rect 37648 27344 37700 27396
rect 37924 27387 37976 27396
rect 37924 27353 37933 27387
rect 37933 27353 37967 27387
rect 37967 27353 37976 27387
rect 37924 27344 37976 27353
rect 38292 27344 38344 27396
rect 29552 27276 29604 27328
rect 30472 27276 30524 27328
rect 31484 27319 31536 27328
rect 31484 27285 31493 27319
rect 31493 27285 31527 27319
rect 31527 27285 31536 27319
rect 31484 27276 31536 27285
rect 33968 27276 34020 27328
rect 35808 27276 35860 27328
rect 38476 27319 38528 27328
rect 38476 27285 38485 27319
rect 38485 27285 38519 27319
rect 38519 27285 38528 27319
rect 38476 27276 38528 27285
rect 38568 27276 38620 27328
rect 39672 27276 39724 27328
rect 39856 27319 39908 27328
rect 39856 27285 39865 27319
rect 39865 27285 39899 27319
rect 39899 27285 39908 27319
rect 39856 27276 39908 27285
rect 41420 27344 41472 27396
rect 40868 27319 40920 27328
rect 40868 27285 40877 27319
rect 40877 27285 40911 27319
rect 40911 27285 40920 27319
rect 40868 27276 40920 27285
rect 41512 27276 41564 27328
rect 41972 27276 42024 27328
rect 42616 27319 42668 27328
rect 42616 27285 42625 27319
rect 42625 27285 42659 27319
rect 42659 27285 42668 27319
rect 42616 27276 42668 27285
rect 46572 27344 46624 27396
rect 46756 27344 46808 27396
rect 50160 27412 50212 27464
rect 46848 27319 46900 27328
rect 46848 27285 46857 27319
rect 46857 27285 46891 27319
rect 46891 27285 46900 27319
rect 46848 27276 46900 27285
rect 48228 27319 48280 27328
rect 48228 27285 48237 27319
rect 48237 27285 48271 27319
rect 48271 27285 48280 27319
rect 48780 27319 48832 27328
rect 48228 27276 48280 27285
rect 48780 27285 48789 27319
rect 48789 27285 48823 27319
rect 48823 27285 48832 27319
rect 48780 27276 48832 27285
rect 50620 27344 50672 27396
rect 52184 27451 52236 27464
rect 52184 27417 52201 27451
rect 52201 27417 52235 27451
rect 52235 27417 52236 27451
rect 52184 27412 52236 27417
rect 50252 27276 50304 27328
rect 54024 27344 54076 27396
rect 57060 27344 57112 27396
rect 57704 27412 57756 27464
rect 58164 27412 58216 27464
rect 58348 27455 58400 27464
rect 58348 27421 58357 27455
rect 58357 27421 58391 27455
rect 58391 27421 58400 27455
rect 58348 27412 58400 27421
rect 58440 27412 58492 27464
rect 59360 27412 59412 27464
rect 60280 27412 60332 27464
rect 61752 27412 61804 27464
rect 62120 27480 62172 27532
rect 63224 27523 63276 27532
rect 63224 27489 63233 27523
rect 63233 27489 63267 27523
rect 63267 27489 63276 27523
rect 63224 27480 63276 27489
rect 63316 27480 63368 27532
rect 63500 27455 63552 27464
rect 63500 27421 63509 27455
rect 63509 27421 63543 27455
rect 63543 27421 63552 27455
rect 63500 27412 63552 27421
rect 64144 27480 64196 27532
rect 64880 27412 64932 27464
rect 65708 27412 65760 27464
rect 68744 27523 68796 27532
rect 68744 27489 68753 27523
rect 68753 27489 68787 27523
rect 68787 27489 68796 27523
rect 69020 27548 69072 27600
rect 70492 27548 70544 27600
rect 74632 27591 74684 27600
rect 74632 27557 74641 27591
rect 74641 27557 74675 27591
rect 74675 27557 74684 27591
rect 74632 27548 74684 27557
rect 75276 27548 75328 27600
rect 79784 27548 79836 27600
rect 81256 27591 81308 27600
rect 81256 27557 81265 27591
rect 81265 27557 81299 27591
rect 81299 27557 81308 27591
rect 81256 27548 81308 27557
rect 81440 27548 81492 27600
rect 82544 27591 82596 27600
rect 82544 27557 82553 27591
rect 82553 27557 82587 27591
rect 82587 27557 82596 27591
rect 82544 27548 82596 27557
rect 85580 27548 85632 27600
rect 87052 27591 87104 27600
rect 87052 27557 87061 27591
rect 87061 27557 87095 27591
rect 87095 27557 87104 27591
rect 87052 27548 87104 27557
rect 87696 27591 87748 27600
rect 87696 27557 87705 27591
rect 87705 27557 87739 27591
rect 87739 27557 87748 27591
rect 87696 27548 87748 27557
rect 68744 27480 68796 27489
rect 70400 27480 70452 27532
rect 65892 27412 65944 27464
rect 66628 27412 66680 27464
rect 69296 27455 69348 27464
rect 69296 27421 69305 27455
rect 69305 27421 69339 27455
rect 69339 27421 69348 27455
rect 69296 27412 69348 27421
rect 69480 27412 69532 27464
rect 70216 27455 70268 27464
rect 70216 27421 70225 27455
rect 70225 27421 70259 27455
rect 70259 27421 70268 27455
rect 71964 27455 72016 27464
rect 70216 27412 70268 27421
rect 58072 27344 58124 27396
rect 50988 27319 51040 27328
rect 50988 27285 50997 27319
rect 50997 27285 51031 27319
rect 51031 27285 51040 27319
rect 50988 27276 51040 27285
rect 51908 27276 51960 27328
rect 53196 27319 53248 27328
rect 53196 27285 53205 27319
rect 53205 27285 53239 27319
rect 53239 27285 53248 27319
rect 53196 27276 53248 27285
rect 53840 27319 53892 27328
rect 53840 27285 53849 27319
rect 53849 27285 53883 27319
rect 53883 27285 53892 27319
rect 53840 27276 53892 27285
rect 55312 27276 55364 27328
rect 55680 27276 55732 27328
rect 56416 27319 56468 27328
rect 56416 27285 56425 27319
rect 56425 27285 56459 27319
rect 56459 27285 56468 27319
rect 56416 27276 56468 27285
rect 57612 27276 57664 27328
rect 59452 27344 59504 27396
rect 59544 27344 59596 27396
rect 59176 27276 59228 27328
rect 60648 27344 60700 27396
rect 60832 27276 60884 27328
rect 62120 27276 62172 27328
rect 64604 27276 64656 27328
rect 66260 27319 66312 27328
rect 66260 27285 66269 27319
rect 66269 27285 66303 27319
rect 66303 27285 66312 27319
rect 66260 27276 66312 27285
rect 68008 27276 68060 27328
rect 68192 27319 68244 27328
rect 68192 27285 68201 27319
rect 68201 27285 68235 27319
rect 68235 27285 68244 27319
rect 68192 27276 68244 27285
rect 68468 27276 68520 27328
rect 69572 27276 69624 27328
rect 71964 27421 71973 27455
rect 71973 27421 72007 27455
rect 72007 27421 72016 27455
rect 71964 27412 72016 27421
rect 72056 27412 72108 27464
rect 72424 27480 72476 27532
rect 74908 27480 74960 27532
rect 75184 27523 75236 27532
rect 75184 27489 75193 27523
rect 75193 27489 75227 27523
rect 75227 27489 75236 27523
rect 75184 27480 75236 27489
rect 75920 27412 75972 27464
rect 76748 27455 76800 27464
rect 76748 27421 76757 27455
rect 76757 27421 76791 27455
rect 76791 27421 76800 27455
rect 76748 27412 76800 27421
rect 76840 27412 76892 27464
rect 78864 27480 78916 27532
rect 79416 27480 79468 27532
rect 84292 27480 84344 27532
rect 85028 27523 85080 27532
rect 70584 27344 70636 27396
rect 78772 27344 78824 27396
rect 79600 27412 79652 27464
rect 80520 27412 80572 27464
rect 81992 27455 82044 27464
rect 81992 27421 82001 27455
rect 82001 27421 82035 27455
rect 82035 27421 82044 27455
rect 81992 27412 82044 27421
rect 82728 27455 82780 27464
rect 82728 27421 82737 27455
rect 82737 27421 82771 27455
rect 82771 27421 82780 27455
rect 82728 27412 82780 27421
rect 83740 27412 83792 27464
rect 83924 27412 83976 27464
rect 85028 27489 85037 27523
rect 85037 27489 85071 27523
rect 85071 27489 85080 27523
rect 85028 27480 85080 27489
rect 85212 27480 85264 27532
rect 90640 27523 90692 27532
rect 90640 27489 90649 27523
rect 90649 27489 90683 27523
rect 90683 27489 90692 27523
rect 90640 27480 90692 27489
rect 91376 27480 91428 27532
rect 94872 27523 94924 27532
rect 70952 27276 71004 27328
rect 71136 27319 71188 27328
rect 71136 27285 71145 27319
rect 71145 27285 71179 27319
rect 71179 27285 71188 27319
rect 71136 27276 71188 27285
rect 71320 27276 71372 27328
rect 74264 27319 74316 27328
rect 74264 27285 74273 27319
rect 74273 27285 74307 27319
rect 74307 27285 74316 27319
rect 74264 27276 74316 27285
rect 74540 27276 74592 27328
rect 74632 27276 74684 27328
rect 76012 27276 76064 27328
rect 78588 27276 78640 27328
rect 78956 27276 79008 27328
rect 79048 27319 79100 27328
rect 79048 27285 79057 27319
rect 79057 27285 79091 27319
rect 79091 27285 79100 27319
rect 79048 27276 79100 27285
rect 79324 27276 79376 27328
rect 84292 27276 84344 27328
rect 84476 27319 84528 27328
rect 84476 27285 84485 27319
rect 84485 27285 84519 27319
rect 84519 27285 84528 27319
rect 84476 27276 84528 27285
rect 86132 27344 86184 27396
rect 86408 27455 86460 27464
rect 86408 27421 86417 27455
rect 86417 27421 86451 27455
rect 86451 27421 86460 27455
rect 87236 27455 87288 27464
rect 86408 27412 86460 27421
rect 87236 27421 87245 27455
rect 87245 27421 87279 27455
rect 87279 27421 87288 27455
rect 87236 27412 87288 27421
rect 87328 27412 87380 27464
rect 88340 27412 88392 27464
rect 86960 27344 87012 27396
rect 88800 27319 88852 27328
rect 88800 27285 88809 27319
rect 88809 27285 88843 27319
rect 88843 27285 88852 27319
rect 88800 27276 88852 27285
rect 89444 27344 89496 27396
rect 89720 27344 89772 27396
rect 91468 27412 91520 27464
rect 94596 27412 94648 27464
rect 94872 27489 94881 27523
rect 94881 27489 94915 27523
rect 94915 27489 94924 27523
rect 94872 27480 94924 27489
rect 95792 27548 95844 27600
rect 95976 27548 96028 27600
rect 96896 27548 96948 27600
rect 101680 27625 101689 27659
rect 101689 27625 101723 27659
rect 101723 27625 101732 27659
rect 101680 27616 101732 27625
rect 98000 27591 98052 27600
rect 98000 27557 98009 27591
rect 98009 27557 98043 27591
rect 98043 27557 98052 27591
rect 98000 27548 98052 27557
rect 98552 27480 98604 27532
rect 99840 27548 99892 27600
rect 100944 27548 100996 27600
rect 103152 27591 103204 27600
rect 103152 27557 103161 27591
rect 103161 27557 103195 27591
rect 103195 27557 103204 27591
rect 103152 27548 103204 27557
rect 105636 27548 105688 27600
rect 107660 27548 107712 27600
rect 109040 27548 109092 27600
rect 113640 27591 113692 27600
rect 113640 27557 113649 27591
rect 113649 27557 113683 27591
rect 113683 27557 113692 27591
rect 113640 27548 113692 27557
rect 115572 27591 115624 27600
rect 115572 27557 115581 27591
rect 115581 27557 115615 27591
rect 115615 27557 115624 27591
rect 115572 27548 115624 27557
rect 92756 27387 92808 27396
rect 90088 27319 90140 27328
rect 90088 27285 90097 27319
rect 90097 27285 90131 27319
rect 90131 27285 90140 27319
rect 90088 27276 90140 27285
rect 90180 27276 90232 27328
rect 92756 27353 92765 27387
rect 92765 27353 92799 27387
rect 92799 27353 92808 27387
rect 92756 27344 92808 27353
rect 96712 27455 96764 27464
rect 96712 27421 96721 27455
rect 96721 27421 96755 27455
rect 96755 27421 96764 27455
rect 96712 27412 96764 27421
rect 91008 27276 91060 27328
rect 91928 27319 91980 27328
rect 91928 27285 91937 27319
rect 91937 27285 91971 27319
rect 91971 27285 91980 27319
rect 91928 27276 91980 27285
rect 92848 27319 92900 27328
rect 92848 27285 92857 27319
rect 92857 27285 92891 27319
rect 92891 27285 92900 27319
rect 92848 27276 92900 27285
rect 94412 27276 94464 27328
rect 94688 27319 94740 27328
rect 94688 27285 94697 27319
rect 94697 27285 94731 27319
rect 94731 27285 94740 27319
rect 94688 27276 94740 27285
rect 94872 27276 94924 27328
rect 96252 27276 96304 27328
rect 96436 27344 96488 27396
rect 98184 27455 98236 27464
rect 98184 27421 98193 27455
rect 98193 27421 98227 27455
rect 98227 27421 98236 27455
rect 98184 27412 98236 27421
rect 99380 27455 99432 27464
rect 99380 27421 99389 27455
rect 99389 27421 99423 27455
rect 99423 27421 99432 27455
rect 99380 27412 99432 27421
rect 99564 27412 99616 27464
rect 101128 27412 101180 27464
rect 102692 27455 102744 27464
rect 102692 27421 102701 27455
rect 102701 27421 102735 27455
rect 102735 27421 102744 27455
rect 102692 27412 102744 27421
rect 102784 27412 102836 27464
rect 105360 27455 105412 27464
rect 105360 27421 105369 27455
rect 105369 27421 105403 27455
rect 105403 27421 105412 27455
rect 105360 27412 105412 27421
rect 106372 27412 106424 27464
rect 106924 27412 106976 27464
rect 97172 27344 97224 27396
rect 100944 27344 100996 27396
rect 104716 27387 104768 27396
rect 104716 27353 104725 27387
rect 104725 27353 104759 27387
rect 104759 27353 104768 27387
rect 104716 27344 104768 27353
rect 104992 27344 105044 27396
rect 110972 27480 111024 27532
rect 116768 27480 116820 27532
rect 108488 27455 108540 27464
rect 108488 27421 108497 27455
rect 108497 27421 108531 27455
rect 108531 27421 108540 27455
rect 108488 27412 108540 27421
rect 109592 27455 109644 27464
rect 109592 27421 109601 27455
rect 109601 27421 109635 27455
rect 109635 27421 109644 27455
rect 109592 27412 109644 27421
rect 109776 27412 109828 27464
rect 111064 27455 111116 27464
rect 111064 27421 111073 27455
rect 111073 27421 111107 27455
rect 111107 27421 111116 27455
rect 111064 27412 111116 27421
rect 112076 27412 112128 27464
rect 114560 27412 114612 27464
rect 116032 27455 116084 27464
rect 116032 27421 116041 27455
rect 116041 27421 116075 27455
rect 116075 27421 116084 27455
rect 116032 27412 116084 27421
rect 117320 27455 117372 27464
rect 117320 27421 117329 27455
rect 117329 27421 117363 27455
rect 117363 27421 117372 27455
rect 117320 27412 117372 27421
rect 96712 27276 96764 27328
rect 104808 27319 104860 27328
rect 104808 27285 104817 27319
rect 104817 27285 104851 27319
rect 104851 27285 104860 27319
rect 104808 27276 104860 27285
rect 104900 27276 104952 27328
rect 105636 27276 105688 27328
rect 110052 27319 110104 27328
rect 110052 27285 110061 27319
rect 110061 27285 110095 27319
rect 110095 27285 110104 27319
rect 110052 27276 110104 27285
rect 112536 27319 112588 27328
rect 112536 27285 112545 27319
rect 112545 27285 112579 27319
rect 112579 27285 112588 27319
rect 112536 27276 112588 27285
rect 114744 27276 114796 27328
rect 115204 27276 115256 27328
rect 30398 27174 30450 27226
rect 30462 27174 30514 27226
rect 30526 27174 30578 27226
rect 30590 27174 30642 27226
rect 30654 27174 30706 27226
rect 59846 27174 59898 27226
rect 59910 27174 59962 27226
rect 59974 27174 60026 27226
rect 60038 27174 60090 27226
rect 60102 27174 60154 27226
rect 89294 27174 89346 27226
rect 89358 27174 89410 27226
rect 89422 27174 89474 27226
rect 89486 27174 89538 27226
rect 89550 27174 89602 27226
rect 1032 27072 1084 27124
rect 4620 27115 4672 27124
rect 4620 27081 4629 27115
rect 4629 27081 4663 27115
rect 4663 27081 4672 27115
rect 4620 27072 4672 27081
rect 7840 27115 7892 27124
rect 7840 27081 7849 27115
rect 7849 27081 7883 27115
rect 7883 27081 7892 27115
rect 7840 27072 7892 27081
rect 9680 27072 9732 27124
rect 11612 27072 11664 27124
rect 1308 26936 1360 26988
rect 2872 26979 2924 26988
rect 2872 26945 2881 26979
rect 2881 26945 2915 26979
rect 2915 26945 2924 26979
rect 2872 26936 2924 26945
rect 3516 26979 3568 26988
rect 3516 26945 3525 26979
rect 3525 26945 3559 26979
rect 3559 26945 3568 26979
rect 3516 26936 3568 26945
rect 4804 26979 4856 26988
rect 4804 26945 4813 26979
rect 4813 26945 4847 26979
rect 4847 26945 4856 26979
rect 4804 26936 4856 26945
rect 1676 26911 1728 26920
rect 1676 26877 1685 26911
rect 1685 26877 1719 26911
rect 1719 26877 1728 26911
rect 1676 26868 1728 26877
rect 10232 26936 10284 26988
rect 26976 27072 27028 27124
rect 29184 27072 29236 27124
rect 11980 27004 12032 27056
rect 14464 27004 14516 27056
rect 15476 27004 15528 27056
rect 17132 27004 17184 27056
rect 19708 27004 19760 27056
rect 22376 27004 22428 27056
rect 26792 27004 26844 27056
rect 27068 27004 27120 27056
rect 29276 27004 29328 27056
rect 14280 26979 14332 26988
rect 14280 26945 14289 26979
rect 14289 26945 14323 26979
rect 14323 26945 14332 26979
rect 14280 26936 14332 26945
rect 19800 26936 19852 26988
rect 20720 26979 20772 26988
rect 20720 26945 20729 26979
rect 20729 26945 20763 26979
rect 20763 26945 20772 26979
rect 20720 26936 20772 26945
rect 27344 26979 27396 26988
rect 27344 26945 27353 26979
rect 27353 26945 27387 26979
rect 27387 26945 27396 26979
rect 27344 26936 27396 26945
rect 30472 27072 30524 27124
rect 32680 27072 32732 27124
rect 32864 27072 32916 27124
rect 33876 27115 33928 27124
rect 33876 27081 33885 27115
rect 33885 27081 33919 27115
rect 33919 27081 33928 27115
rect 33876 27072 33928 27081
rect 31852 27004 31904 27056
rect 33968 27004 34020 27056
rect 29552 26979 29604 26988
rect 24124 26868 24176 26920
rect 27160 26868 27212 26920
rect 29552 26945 29561 26979
rect 29561 26945 29595 26979
rect 29595 26945 29604 26979
rect 29552 26936 29604 26945
rect 27528 26868 27580 26920
rect 29000 26868 29052 26920
rect 29368 26868 29420 26920
rect 30748 26936 30800 26988
rect 32036 26936 32088 26988
rect 32128 26936 32180 26988
rect 35440 27072 35492 27124
rect 38108 27115 38160 27124
rect 38108 27081 38117 27115
rect 38117 27081 38151 27115
rect 38151 27081 38160 27115
rect 38108 27072 38160 27081
rect 38200 27072 38252 27124
rect 40316 27072 40368 27124
rect 40500 27115 40552 27124
rect 40500 27081 40509 27115
rect 40509 27081 40543 27115
rect 40543 27081 40552 27115
rect 40500 27072 40552 27081
rect 41328 27115 41380 27124
rect 41328 27081 41337 27115
rect 41337 27081 41371 27115
rect 41371 27081 41380 27115
rect 41328 27072 41380 27081
rect 41604 27072 41656 27124
rect 45652 27072 45704 27124
rect 45836 27115 45888 27124
rect 45836 27081 45845 27115
rect 45845 27081 45879 27115
rect 45879 27081 45888 27115
rect 45836 27072 45888 27081
rect 52920 27115 52972 27124
rect 34888 27004 34940 27056
rect 34612 26979 34664 26988
rect 34612 26945 34621 26979
rect 34621 26945 34655 26979
rect 34655 26945 34664 26979
rect 34612 26936 34664 26945
rect 35716 26979 35768 26988
rect 35716 26945 35725 26979
rect 35725 26945 35759 26979
rect 35759 26945 35768 26979
rect 35716 26936 35768 26945
rect 35808 26936 35860 26988
rect 36636 26979 36688 26988
rect 36636 26945 36645 26979
rect 36645 26945 36679 26979
rect 36679 26945 36688 26979
rect 36636 26936 36688 26945
rect 41880 27004 41932 27056
rect 38384 26936 38436 26988
rect 2964 26800 3016 26852
rect 9404 26800 9456 26852
rect 10508 26800 10560 26852
rect 9588 26732 9640 26784
rect 15568 26732 15620 26784
rect 16028 26800 16080 26852
rect 17040 26800 17092 26852
rect 20536 26843 20588 26852
rect 20536 26809 20545 26843
rect 20545 26809 20579 26843
rect 20579 26809 20588 26843
rect 20536 26800 20588 26809
rect 22008 26800 22060 26852
rect 22192 26800 22244 26852
rect 22284 26800 22336 26852
rect 26792 26800 26844 26852
rect 27252 26800 27304 26852
rect 29092 26800 29144 26852
rect 29552 26800 29604 26852
rect 33600 26800 33652 26852
rect 21088 26732 21140 26784
rect 21916 26732 21968 26784
rect 27068 26732 27120 26784
rect 27160 26732 27212 26784
rect 29276 26732 29328 26784
rect 30104 26732 30156 26784
rect 34060 26732 34112 26784
rect 34980 26800 35032 26852
rect 39304 26868 39356 26920
rect 39856 26936 39908 26988
rect 41420 26936 41472 26988
rect 46480 27004 46532 27056
rect 46572 27004 46624 27056
rect 46848 27004 46900 27056
rect 50620 27004 50672 27056
rect 50712 27047 50764 27056
rect 50712 27013 50721 27047
rect 50721 27013 50755 27047
rect 50755 27013 50764 27047
rect 50712 27004 50764 27013
rect 51172 27004 51224 27056
rect 39672 26868 39724 26920
rect 41236 26868 41288 26920
rect 46204 26936 46256 26988
rect 41696 26868 41748 26920
rect 48504 26868 48556 26920
rect 48964 26936 49016 26988
rect 50068 26936 50120 26988
rect 50344 26936 50396 26988
rect 50712 26868 50764 26920
rect 44088 26800 44140 26852
rect 45928 26800 45980 26852
rect 49976 26843 50028 26852
rect 46940 26775 46992 26784
rect 46940 26741 46949 26775
rect 46949 26741 46983 26775
rect 46983 26741 46992 26775
rect 46940 26732 46992 26741
rect 47124 26732 47176 26784
rect 49056 26732 49108 26784
rect 49148 26732 49200 26784
rect 49976 26809 49985 26843
rect 49985 26809 50019 26843
rect 50019 26809 50028 26843
rect 49976 26800 50028 26809
rect 50160 26800 50212 26852
rect 51724 26868 51776 26920
rect 52920 27081 52929 27115
rect 52929 27081 52963 27115
rect 52963 27081 52972 27115
rect 52920 27072 52972 27081
rect 53012 27072 53064 27124
rect 53288 27004 53340 27056
rect 53840 27004 53892 27056
rect 54024 27072 54076 27124
rect 55404 27072 55456 27124
rect 56508 27115 56560 27124
rect 56508 27081 56517 27115
rect 56517 27081 56551 27115
rect 56551 27081 56560 27115
rect 56508 27072 56560 27081
rect 57520 27072 57572 27124
rect 58072 27072 58124 27124
rect 58532 27072 58584 27124
rect 59176 27115 59228 27124
rect 59176 27081 59185 27115
rect 59185 27081 59219 27115
rect 59219 27081 59228 27115
rect 59176 27072 59228 27081
rect 59084 27004 59136 27056
rect 59452 27004 59504 27056
rect 70492 27072 70544 27124
rect 71136 27072 71188 27124
rect 74540 27072 74592 27124
rect 74724 27072 74776 27124
rect 62948 27004 63000 27056
rect 53932 26911 53984 26920
rect 53932 26877 53941 26911
rect 53941 26877 53975 26911
rect 53975 26877 53984 26911
rect 53932 26868 53984 26877
rect 51632 26732 51684 26784
rect 54024 26800 54076 26852
rect 55128 26936 55180 26988
rect 55496 26936 55548 26988
rect 55680 26979 55732 26988
rect 55680 26945 55689 26979
rect 55689 26945 55723 26979
rect 55723 26945 55732 26979
rect 55680 26936 55732 26945
rect 56324 26979 56376 26988
rect 56324 26945 56333 26979
rect 56333 26945 56367 26979
rect 56367 26945 56376 26979
rect 56324 26936 56376 26945
rect 56692 26979 56744 26988
rect 56692 26945 56701 26979
rect 56701 26945 56735 26979
rect 56735 26945 56744 26979
rect 56692 26936 56744 26945
rect 57336 26979 57388 26988
rect 57336 26945 57345 26979
rect 57345 26945 57379 26979
rect 57379 26945 57388 26979
rect 57336 26936 57388 26945
rect 54300 26868 54352 26920
rect 55864 26911 55916 26920
rect 55864 26877 55873 26911
rect 55873 26877 55907 26911
rect 55907 26877 55916 26911
rect 55864 26868 55916 26877
rect 57244 26868 57296 26920
rect 59176 26936 59228 26988
rect 59360 26936 59412 26988
rect 58072 26868 58124 26920
rect 58256 26868 58308 26920
rect 59636 26936 59688 26988
rect 60188 26936 60240 26988
rect 58164 26843 58216 26852
rect 58164 26809 58173 26843
rect 58173 26809 58207 26843
rect 58207 26809 58216 26843
rect 58164 26800 58216 26809
rect 59544 26868 59596 26920
rect 61752 26936 61804 26988
rect 61936 26979 61988 26988
rect 61936 26945 61945 26979
rect 61945 26945 61979 26979
rect 61979 26945 61988 26979
rect 61936 26936 61988 26945
rect 62580 26979 62632 26988
rect 62580 26945 62589 26979
rect 62589 26945 62623 26979
rect 62623 26945 62632 26979
rect 63684 26979 63736 26988
rect 62580 26936 62632 26945
rect 63684 26945 63693 26979
rect 63693 26945 63727 26979
rect 63727 26945 63736 26979
rect 63684 26936 63736 26945
rect 64604 26936 64656 26988
rect 64696 26936 64748 26988
rect 60464 26868 60516 26920
rect 62212 26911 62264 26920
rect 62212 26877 62221 26911
rect 62221 26877 62255 26911
rect 62255 26877 62264 26911
rect 62212 26868 62264 26877
rect 62396 26868 62448 26920
rect 60556 26800 60608 26852
rect 54300 26732 54352 26784
rect 54392 26732 54444 26784
rect 60648 26732 60700 26784
rect 61200 26800 61252 26852
rect 64696 26800 64748 26852
rect 64880 26868 64932 26920
rect 61476 26732 61528 26784
rect 61844 26732 61896 26784
rect 61936 26732 61988 26784
rect 63224 26732 63276 26784
rect 64052 26732 64104 26784
rect 64144 26732 64196 26784
rect 65984 26936 66036 26988
rect 68192 27004 68244 27056
rect 71872 27004 71924 27056
rect 68836 26936 68888 26988
rect 69112 26936 69164 26988
rect 69848 26868 69900 26920
rect 70676 26936 70728 26988
rect 70952 26979 71004 26988
rect 70952 26945 70961 26979
rect 70961 26945 70995 26979
rect 70995 26945 71004 26979
rect 70952 26936 71004 26945
rect 72608 26936 72660 26988
rect 73160 26979 73212 26988
rect 73160 26945 73169 26979
rect 73169 26945 73203 26979
rect 73203 26945 73212 26979
rect 73160 26936 73212 26945
rect 74448 26936 74500 26988
rect 75000 27004 75052 27056
rect 76564 27004 76616 27056
rect 77300 27072 77352 27124
rect 74816 26936 74868 26988
rect 79232 27072 79284 27124
rect 79876 27072 79928 27124
rect 83924 27072 83976 27124
rect 84200 27072 84252 27124
rect 84936 27072 84988 27124
rect 89076 27072 89128 27124
rect 85672 27004 85724 27056
rect 79048 26936 79100 26988
rect 70308 26800 70360 26852
rect 71872 26843 71924 26852
rect 71872 26809 71881 26843
rect 71881 26809 71915 26843
rect 71915 26809 71924 26843
rect 71872 26800 71924 26809
rect 75920 26868 75972 26920
rect 76104 26911 76156 26920
rect 76104 26877 76113 26911
rect 76113 26877 76147 26911
rect 76147 26877 76156 26911
rect 76104 26868 76156 26877
rect 76196 26911 76248 26920
rect 76196 26877 76205 26911
rect 76205 26877 76239 26911
rect 76239 26877 76248 26911
rect 76196 26868 76248 26877
rect 80060 26936 80112 26988
rect 84016 26936 84068 26988
rect 78680 26800 78732 26852
rect 84844 26868 84896 26920
rect 66260 26732 66312 26784
rect 69112 26732 69164 26784
rect 69572 26732 69624 26784
rect 70400 26732 70452 26784
rect 70768 26775 70820 26784
rect 70768 26741 70777 26775
rect 70777 26741 70811 26775
rect 70811 26741 70820 26775
rect 70768 26732 70820 26741
rect 72516 26732 72568 26784
rect 72700 26732 72752 26784
rect 73068 26732 73120 26784
rect 75552 26732 75604 26784
rect 76472 26732 76524 26784
rect 76564 26732 76616 26784
rect 78404 26732 78456 26784
rect 84568 26800 84620 26852
rect 79508 26732 79560 26784
rect 85304 26936 85356 26988
rect 86960 27004 87012 27056
rect 90088 27004 90140 27056
rect 90732 27072 90784 27124
rect 92480 27072 92532 27124
rect 95240 27072 95292 27124
rect 95792 27072 95844 27124
rect 99564 27072 99616 27124
rect 100576 27115 100628 27124
rect 100576 27081 100585 27115
rect 100585 27081 100619 27115
rect 100619 27081 100628 27115
rect 100576 27072 100628 27081
rect 104624 27072 104676 27124
rect 94412 27047 94464 27056
rect 85212 26868 85264 26920
rect 89168 26936 89220 26988
rect 89628 26979 89680 26988
rect 89628 26945 89637 26979
rect 89637 26945 89671 26979
rect 89671 26945 89680 26979
rect 89628 26936 89680 26945
rect 90180 26936 90232 26988
rect 90364 26936 90416 26988
rect 90640 26936 90692 26988
rect 91376 26979 91428 26988
rect 91376 26945 91385 26979
rect 91385 26945 91419 26979
rect 91419 26945 91428 26979
rect 91376 26936 91428 26945
rect 94412 27013 94421 27047
rect 94421 27013 94455 27047
rect 94455 27013 94464 27047
rect 94412 27004 94464 27013
rect 94596 27004 94648 27056
rect 101680 27004 101732 27056
rect 104716 27047 104768 27056
rect 104716 27013 104725 27047
rect 104725 27013 104759 27047
rect 104759 27013 104768 27047
rect 110052 27072 110104 27124
rect 111524 27115 111576 27124
rect 111524 27081 111533 27115
rect 111533 27081 111567 27115
rect 111567 27081 111576 27115
rect 111524 27072 111576 27081
rect 117228 27072 117280 27124
rect 116768 27047 116820 27056
rect 104716 27004 104768 27013
rect 116768 27013 116777 27047
rect 116777 27013 116811 27047
rect 116811 27013 116820 27047
rect 116768 27004 116820 27013
rect 94872 26936 94924 26988
rect 95240 26979 95292 26988
rect 95240 26945 95249 26979
rect 95249 26945 95283 26979
rect 95283 26945 95292 26979
rect 95240 26936 95292 26945
rect 95884 26979 95936 26988
rect 95884 26945 95893 26979
rect 95893 26945 95927 26979
rect 95927 26945 95936 26979
rect 95884 26936 95936 26945
rect 95976 26936 96028 26988
rect 86132 26800 86184 26852
rect 91744 26868 91796 26920
rect 100852 26936 100904 26988
rect 103336 26936 103388 26988
rect 105544 26979 105596 26988
rect 105544 26945 105553 26979
rect 105553 26945 105587 26979
rect 105587 26945 105596 26979
rect 105544 26936 105596 26945
rect 111708 26979 111760 26988
rect 111708 26945 111717 26979
rect 111717 26945 111751 26979
rect 111751 26945 111760 26979
rect 111708 26936 111760 26945
rect 91836 26800 91888 26852
rect 92204 26843 92256 26852
rect 92204 26809 92213 26843
rect 92213 26809 92247 26843
rect 92247 26809 92256 26843
rect 92204 26800 92256 26809
rect 94044 26800 94096 26852
rect 85396 26775 85448 26784
rect 85396 26741 85405 26775
rect 85405 26741 85439 26775
rect 85439 26741 85448 26775
rect 85396 26732 85448 26741
rect 86224 26732 86276 26784
rect 86868 26732 86920 26784
rect 90088 26732 90140 26784
rect 90732 26732 90784 26784
rect 90916 26775 90968 26784
rect 90916 26741 90925 26775
rect 90925 26741 90959 26775
rect 90959 26741 90968 26775
rect 90916 26732 90968 26741
rect 91744 26732 91796 26784
rect 100208 26800 100260 26852
rect 104348 26868 104400 26920
rect 108488 26868 108540 26920
rect 109592 26868 109644 26920
rect 113640 26868 113692 26920
rect 104900 26843 104952 26852
rect 104900 26809 104909 26843
rect 104909 26809 104943 26843
rect 104943 26809 104952 26843
rect 104900 26800 104952 26809
rect 117136 26936 117188 26988
rect 117964 26979 118016 26988
rect 117964 26945 117973 26979
rect 117973 26945 118007 26979
rect 118007 26945 118016 26979
rect 117964 26936 118016 26945
rect 117780 26732 117832 26784
rect 15674 26630 15726 26682
rect 15738 26630 15790 26682
rect 15802 26630 15854 26682
rect 15866 26630 15918 26682
rect 15930 26630 15982 26682
rect 45122 26630 45174 26682
rect 45186 26630 45238 26682
rect 45250 26630 45302 26682
rect 45314 26630 45366 26682
rect 45378 26630 45430 26682
rect 74570 26630 74622 26682
rect 74634 26630 74686 26682
rect 74698 26630 74750 26682
rect 74762 26630 74814 26682
rect 74826 26630 74878 26682
rect 104018 26630 104070 26682
rect 104082 26630 104134 26682
rect 104146 26630 104198 26682
rect 104210 26630 104262 26682
rect 104274 26630 104326 26682
rect 1676 26528 1728 26580
rect 22100 26528 22152 26580
rect 24124 26528 24176 26580
rect 29552 26528 29604 26580
rect 29736 26571 29788 26580
rect 29736 26537 29745 26571
rect 29745 26537 29779 26571
rect 29779 26537 29788 26571
rect 29736 26528 29788 26537
rect 31484 26528 31536 26580
rect 40960 26528 41012 26580
rect 41236 26528 41288 26580
rect 46204 26528 46256 26580
rect 46572 26528 46624 26580
rect 46756 26528 46808 26580
rect 50896 26528 50948 26580
rect 51172 26528 51224 26580
rect 60556 26528 60608 26580
rect 61752 26528 61804 26580
rect 68376 26528 68428 26580
rect 68468 26528 68520 26580
rect 70032 26571 70084 26580
rect 70032 26537 70041 26571
rect 70041 26537 70075 26571
rect 70075 26537 70084 26571
rect 70032 26528 70084 26537
rect 2780 26460 2832 26512
rect 15568 26460 15620 26512
rect 21180 26460 21232 26512
rect 22376 26460 22428 26512
rect 30104 26460 30156 26512
rect 30196 26460 30248 26512
rect 31760 26460 31812 26512
rect 31852 26460 31904 26512
rect 43444 26460 43496 26512
rect 45652 26460 45704 26512
rect 48228 26460 48280 26512
rect 50804 26460 50856 26512
rect 1216 26392 1268 26444
rect 6644 26392 6696 26444
rect 24124 26392 24176 26444
rect 28172 26392 28224 26444
rect 31576 26392 31628 26444
rect 31668 26392 31720 26444
rect 35808 26435 35860 26444
rect 22376 26324 22428 26376
rect 20 26188 72 26240
rect 2872 26188 2924 26240
rect 9036 26188 9088 26240
rect 10324 26188 10376 26240
rect 29460 26324 29512 26376
rect 29644 26324 29696 26376
rect 24492 26256 24544 26308
rect 35532 26324 35584 26376
rect 35808 26401 35817 26435
rect 35817 26401 35851 26435
rect 35851 26401 35860 26435
rect 35808 26392 35860 26401
rect 35900 26392 35952 26444
rect 40776 26392 40828 26444
rect 41236 26392 41288 26444
rect 41052 26324 41104 26376
rect 51448 26460 51500 26512
rect 54760 26460 54812 26512
rect 56324 26460 56376 26512
rect 57336 26460 57388 26512
rect 58716 26503 58768 26512
rect 58716 26469 58725 26503
rect 58725 26469 58759 26503
rect 58759 26469 58768 26503
rect 58716 26460 58768 26469
rect 54392 26392 54444 26444
rect 70492 26460 70544 26512
rect 74724 26460 74776 26512
rect 74908 26528 74960 26580
rect 76564 26528 76616 26580
rect 77392 26571 77444 26580
rect 77392 26537 77401 26571
rect 77401 26537 77435 26571
rect 77435 26537 77444 26571
rect 77392 26528 77444 26537
rect 78404 26528 78456 26580
rect 79508 26528 79560 26580
rect 46664 26367 46716 26376
rect 46664 26333 46673 26367
rect 46673 26333 46707 26367
rect 46707 26333 46716 26367
rect 46664 26324 46716 26333
rect 48228 26367 48280 26376
rect 48228 26333 48237 26367
rect 48237 26333 48271 26367
rect 48271 26333 48280 26367
rect 48228 26324 48280 26333
rect 49240 26367 49292 26376
rect 49240 26333 49249 26367
rect 49249 26333 49283 26367
rect 49283 26333 49292 26367
rect 49240 26324 49292 26333
rect 50344 26367 50396 26376
rect 50344 26333 50353 26367
rect 50353 26333 50387 26367
rect 50387 26333 50396 26367
rect 53748 26367 53800 26376
rect 50344 26324 50396 26333
rect 53748 26333 53757 26367
rect 53757 26333 53791 26367
rect 53791 26333 53800 26367
rect 53748 26324 53800 26333
rect 61752 26392 61804 26444
rect 30104 26256 30156 26308
rect 31760 26256 31812 26308
rect 26792 26188 26844 26240
rect 35716 26256 35768 26308
rect 40960 26256 41012 26308
rect 41420 26256 41472 26308
rect 46848 26256 46900 26308
rect 47308 26256 47360 26308
rect 50988 26256 51040 26308
rect 51264 26256 51316 26308
rect 53380 26256 53432 26308
rect 53564 26256 53616 26308
rect 56876 26324 56928 26376
rect 61016 26324 61068 26376
rect 61108 26324 61160 26376
rect 35164 26231 35216 26240
rect 35164 26197 35173 26231
rect 35173 26197 35207 26231
rect 35207 26197 35216 26231
rect 35164 26188 35216 26197
rect 35348 26188 35400 26240
rect 37648 26188 37700 26240
rect 40224 26188 40276 26240
rect 49976 26188 50028 26240
rect 50160 26231 50212 26240
rect 50160 26197 50169 26231
rect 50169 26197 50203 26231
rect 50203 26197 50212 26231
rect 50160 26188 50212 26197
rect 50528 26188 50580 26240
rect 59176 26256 59228 26308
rect 60740 26256 60792 26308
rect 55680 26188 55732 26240
rect 60464 26188 60516 26240
rect 60556 26188 60608 26240
rect 61936 26256 61988 26308
rect 63500 26392 63552 26444
rect 69940 26392 69992 26444
rect 68560 26324 68612 26376
rect 68652 26324 68704 26376
rect 70768 26324 70820 26376
rect 71780 26324 71832 26376
rect 72240 26392 72292 26444
rect 77484 26392 77536 26444
rect 79048 26460 79100 26512
rect 84016 26528 84068 26580
rect 85304 26528 85356 26580
rect 85396 26528 85448 26580
rect 100852 26528 100904 26580
rect 104348 26528 104400 26580
rect 110972 26528 111024 26580
rect 90088 26460 90140 26512
rect 74908 26324 74960 26376
rect 75092 26324 75144 26376
rect 76472 26367 76524 26376
rect 76472 26333 76481 26367
rect 76481 26333 76515 26367
rect 76515 26333 76524 26367
rect 76472 26324 76524 26333
rect 77576 26367 77628 26376
rect 77576 26333 77585 26367
rect 77585 26333 77619 26367
rect 77619 26333 77628 26367
rect 77576 26324 77628 26333
rect 78680 26324 78732 26376
rect 70676 26188 70728 26240
rect 71320 26256 71372 26308
rect 71596 26256 71648 26308
rect 72792 26256 72844 26308
rect 79692 26324 79744 26376
rect 82268 26392 82320 26444
rect 81900 26324 81952 26376
rect 89076 26324 89128 26376
rect 71044 26188 71096 26240
rect 71780 26188 71832 26240
rect 71872 26231 71924 26240
rect 71872 26197 71881 26231
rect 71881 26197 71915 26231
rect 71915 26197 71924 26231
rect 71872 26188 71924 26197
rect 74724 26188 74776 26240
rect 76656 26231 76708 26240
rect 76656 26197 76665 26231
rect 76665 26197 76699 26231
rect 76699 26197 76708 26231
rect 76656 26188 76708 26197
rect 79600 26231 79652 26240
rect 79600 26197 79609 26231
rect 79609 26197 79643 26231
rect 79643 26197 79652 26231
rect 79600 26188 79652 26197
rect 81164 26256 81216 26308
rect 89168 26256 89220 26308
rect 89996 26324 90048 26376
rect 90180 26392 90232 26444
rect 91744 26392 91796 26444
rect 95792 26460 95844 26512
rect 103336 26460 103388 26512
rect 117412 26460 117464 26512
rect 90456 26367 90508 26376
rect 90456 26333 90465 26367
rect 90465 26333 90499 26367
rect 90499 26333 90508 26367
rect 93676 26367 93728 26376
rect 90456 26324 90508 26333
rect 89352 26256 89404 26308
rect 90272 26231 90324 26240
rect 90272 26197 90281 26231
rect 90281 26197 90315 26231
rect 90315 26197 90324 26231
rect 90272 26188 90324 26197
rect 91836 26299 91888 26308
rect 91836 26265 91845 26299
rect 91845 26265 91879 26299
rect 91879 26265 91888 26299
rect 93676 26333 93685 26367
rect 93685 26333 93719 26367
rect 93719 26333 93728 26367
rect 93676 26324 93728 26333
rect 102784 26392 102836 26444
rect 116860 26324 116912 26376
rect 117044 26324 117096 26376
rect 118516 26324 118568 26376
rect 91836 26256 91888 26265
rect 117780 26256 117832 26308
rect 118056 26256 118108 26308
rect 93492 26231 93544 26240
rect 93492 26197 93501 26231
rect 93501 26197 93535 26231
rect 93535 26197 93544 26231
rect 93492 26188 93544 26197
rect 30398 26086 30450 26138
rect 30462 26086 30514 26138
rect 30526 26086 30578 26138
rect 30590 26086 30642 26138
rect 30654 26086 30706 26138
rect 59846 26086 59898 26138
rect 59910 26086 59962 26138
rect 59974 26086 60026 26138
rect 60038 26086 60090 26138
rect 60102 26086 60154 26138
rect 89294 26086 89346 26138
rect 89358 26086 89410 26138
rect 89422 26086 89474 26138
rect 89486 26086 89538 26138
rect 89550 26086 89602 26138
rect 1400 26027 1452 26036
rect 1400 25993 1409 26027
rect 1409 25993 1443 26027
rect 1443 25993 1452 26027
rect 1400 25984 1452 25993
rect 29092 25984 29144 26036
rect 31668 25984 31720 26036
rect 31760 25984 31812 26036
rect 34888 25984 34940 26036
rect 36636 25984 36688 26036
rect 50804 25984 50856 26036
rect 55680 25984 55732 26036
rect 60280 25984 60332 26036
rect 63316 25984 63368 26036
rect 68560 25984 68612 26036
rect 72056 25984 72108 26036
rect 76104 26027 76156 26036
rect 76104 25993 76113 26027
rect 76113 25993 76147 26027
rect 76147 25993 76156 26027
rect 76104 25984 76156 25993
rect 77484 25984 77536 26036
rect 85028 25984 85080 26036
rect 54484 25916 54536 25968
rect 35256 25848 35308 25900
rect 40960 25848 41012 25900
rect 46756 25848 46808 25900
rect 49976 25848 50028 25900
rect 54116 25848 54168 25900
rect 58164 25916 58216 25968
rect 68284 25916 68336 25968
rect 71320 25916 71372 25968
rect 81164 25916 81216 25968
rect 58072 25891 58124 25900
rect 58072 25857 58081 25891
rect 58081 25857 58115 25891
rect 58115 25857 58124 25891
rect 58072 25848 58124 25857
rect 58532 25848 58584 25900
rect 61844 25891 61896 25900
rect 56784 25780 56836 25832
rect 61844 25857 61853 25891
rect 61853 25857 61887 25891
rect 61887 25857 61896 25891
rect 61844 25848 61896 25857
rect 68008 25848 68060 25900
rect 72792 25848 72844 25900
rect 76288 25891 76340 25900
rect 76288 25857 76297 25891
rect 76297 25857 76331 25891
rect 76331 25857 76340 25891
rect 76288 25848 76340 25857
rect 77576 25848 77628 25900
rect 82268 25848 82320 25900
rect 60372 25823 60424 25832
rect 60372 25789 60381 25823
rect 60381 25789 60415 25823
rect 60415 25789 60424 25823
rect 60372 25780 60424 25789
rect 64144 25780 64196 25832
rect 60924 25712 60976 25764
rect 61016 25712 61068 25764
rect 76840 25780 76892 25832
rect 94688 25712 94740 25764
rect 119804 25916 119856 25968
rect 117872 25848 117924 25900
rect 57888 25644 57940 25696
rect 58532 25687 58584 25696
rect 58532 25653 58541 25687
rect 58541 25653 58575 25687
rect 58575 25653 58584 25687
rect 58532 25644 58584 25653
rect 59452 25644 59504 25696
rect 60372 25644 60424 25696
rect 78864 25644 78916 25696
rect 15674 25542 15726 25594
rect 15738 25542 15790 25594
rect 15802 25542 15854 25594
rect 15866 25542 15918 25594
rect 15930 25542 15982 25594
rect 45122 25542 45174 25594
rect 45186 25542 45238 25594
rect 45250 25542 45302 25594
rect 45314 25542 45366 25594
rect 45378 25542 45430 25594
rect 74570 25542 74622 25594
rect 74634 25542 74686 25594
rect 74698 25542 74750 25594
rect 74762 25542 74814 25594
rect 74826 25542 74878 25594
rect 104018 25542 104070 25594
rect 104082 25542 104134 25594
rect 104146 25542 104198 25594
rect 104210 25542 104262 25594
rect 104274 25542 104326 25594
rect 4436 25440 4488 25492
rect 59452 25440 59504 25492
rect 47216 25304 47268 25356
rect 54484 25372 54536 25424
rect 56876 25304 56928 25356
rect 32864 25279 32916 25288
rect 32864 25245 32873 25279
rect 32873 25245 32907 25279
rect 32907 25245 32916 25279
rect 32864 25236 32916 25245
rect 42708 25236 42760 25288
rect 57888 25279 57940 25288
rect 57888 25245 57897 25279
rect 57897 25245 57931 25279
rect 57931 25245 57940 25279
rect 57888 25236 57940 25245
rect 64052 25279 64104 25288
rect 64052 25245 64061 25279
rect 64061 25245 64095 25279
rect 64095 25245 64104 25279
rect 64052 25236 64104 25245
rect 107660 25236 107712 25288
rect 34520 25168 34572 25220
rect 64236 25211 64288 25220
rect 64236 25177 64245 25211
rect 64245 25177 64279 25211
rect 64279 25177 64288 25211
rect 64236 25168 64288 25177
rect 86408 25100 86460 25152
rect 117964 25143 118016 25152
rect 117964 25109 117973 25143
rect 117973 25109 118007 25143
rect 118007 25109 118016 25143
rect 117964 25100 118016 25109
rect 30398 24998 30450 25050
rect 30462 24998 30514 25050
rect 30526 24998 30578 25050
rect 30590 24998 30642 25050
rect 30654 24998 30706 25050
rect 59846 24998 59898 25050
rect 59910 24998 59962 25050
rect 59974 24998 60026 25050
rect 60038 24998 60090 25050
rect 60102 24998 60154 25050
rect 89294 24998 89346 25050
rect 89358 24998 89410 25050
rect 89422 24998 89474 25050
rect 89486 24998 89538 25050
rect 89550 24998 89602 25050
rect 29552 24896 29604 24948
rect 32864 24896 32916 24948
rect 1400 24735 1452 24744
rect 1400 24701 1409 24735
rect 1409 24701 1443 24735
rect 1443 24701 1452 24735
rect 1400 24692 1452 24701
rect 31116 24735 31168 24744
rect 31116 24701 31125 24735
rect 31125 24701 31159 24735
rect 31159 24701 31168 24735
rect 31116 24692 31168 24701
rect 31300 24735 31352 24744
rect 31300 24701 31309 24735
rect 31309 24701 31343 24735
rect 31343 24701 31352 24735
rect 31300 24692 31352 24701
rect 31760 24760 31812 24812
rect 32864 24692 32916 24744
rect 42708 24624 42760 24676
rect 31760 24599 31812 24608
rect 31760 24565 31769 24599
rect 31769 24565 31803 24599
rect 31803 24565 31812 24599
rect 31760 24556 31812 24565
rect 59636 24556 59688 24608
rect 64236 24556 64288 24608
rect 117964 24599 118016 24608
rect 117964 24565 117973 24599
rect 117973 24565 118007 24599
rect 118007 24565 118016 24599
rect 117964 24556 118016 24565
rect 15674 24454 15726 24506
rect 15738 24454 15790 24506
rect 15802 24454 15854 24506
rect 15866 24454 15918 24506
rect 15930 24454 15982 24506
rect 45122 24454 45174 24506
rect 45186 24454 45238 24506
rect 45250 24454 45302 24506
rect 45314 24454 45366 24506
rect 45378 24454 45430 24506
rect 74570 24454 74622 24506
rect 74634 24454 74686 24506
rect 74698 24454 74750 24506
rect 74762 24454 74814 24506
rect 74826 24454 74878 24506
rect 104018 24454 104070 24506
rect 104082 24454 104134 24506
rect 104146 24454 104198 24506
rect 104210 24454 104262 24506
rect 104274 24454 104326 24506
rect 34520 24352 34572 24404
rect 31300 24259 31352 24268
rect 31300 24225 31309 24259
rect 31309 24225 31343 24259
rect 31343 24225 31352 24259
rect 31300 24216 31352 24225
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 1676 24191 1728 24200
rect 1676 24157 1685 24191
rect 1685 24157 1719 24191
rect 1719 24157 1728 24191
rect 1676 24148 1728 24157
rect 2688 24148 2740 24200
rect 2964 24148 3016 24200
rect 51080 24148 51132 24200
rect 51448 24148 51500 24200
rect 35440 24080 35492 24132
rect 102232 24080 102284 24132
rect 1492 24012 1544 24064
rect 28816 24012 28868 24064
rect 30398 23910 30450 23962
rect 30462 23910 30514 23962
rect 30526 23910 30578 23962
rect 30590 23910 30642 23962
rect 30654 23910 30706 23962
rect 59846 23910 59898 23962
rect 59910 23910 59962 23962
rect 59974 23910 60026 23962
rect 60038 23910 60090 23962
rect 60102 23910 60154 23962
rect 89294 23910 89346 23962
rect 89358 23910 89410 23962
rect 89422 23910 89474 23962
rect 89486 23910 89538 23962
rect 89550 23910 89602 23962
rect 1768 23672 1820 23724
rect 91008 23672 91060 23724
rect 117228 23604 117280 23656
rect 1400 23511 1452 23520
rect 1400 23477 1409 23511
rect 1409 23477 1443 23511
rect 1443 23477 1452 23511
rect 1400 23468 1452 23477
rect 15674 23366 15726 23418
rect 15738 23366 15790 23418
rect 15802 23366 15854 23418
rect 15866 23366 15918 23418
rect 15930 23366 15982 23418
rect 45122 23366 45174 23418
rect 45186 23366 45238 23418
rect 45250 23366 45302 23418
rect 45314 23366 45366 23418
rect 45378 23366 45430 23418
rect 74570 23366 74622 23418
rect 74634 23366 74686 23418
rect 74698 23366 74750 23418
rect 74762 23366 74814 23418
rect 74826 23366 74878 23418
rect 104018 23366 104070 23418
rect 104082 23366 104134 23418
rect 104146 23366 104198 23418
rect 104210 23366 104262 23418
rect 104274 23366 104326 23418
rect 1676 22924 1728 22976
rect 11704 22924 11756 22976
rect 14648 22924 14700 22976
rect 71228 22924 71280 22976
rect 30398 22822 30450 22874
rect 30462 22822 30514 22874
rect 30526 22822 30578 22874
rect 30590 22822 30642 22874
rect 30654 22822 30706 22874
rect 59846 22822 59898 22874
rect 59910 22822 59962 22874
rect 59974 22822 60026 22874
rect 60038 22822 60090 22874
rect 60102 22822 60154 22874
rect 89294 22822 89346 22874
rect 89358 22822 89410 22874
rect 89422 22822 89474 22874
rect 89486 22822 89538 22874
rect 89550 22822 89602 22874
rect 9220 22720 9272 22772
rect 98184 22720 98236 22772
rect 88800 22652 88852 22704
rect 94780 22627 94832 22636
rect 94780 22593 94789 22627
rect 94789 22593 94823 22627
rect 94823 22593 94832 22627
rect 94780 22584 94832 22593
rect 94964 22559 95016 22568
rect 94964 22525 94973 22559
rect 94973 22525 95007 22559
rect 95007 22525 95016 22559
rect 94964 22516 95016 22525
rect 117964 22491 118016 22500
rect 117964 22457 117973 22491
rect 117973 22457 118007 22491
rect 118007 22457 118016 22491
rect 117964 22448 118016 22457
rect 15674 22278 15726 22330
rect 15738 22278 15790 22330
rect 15802 22278 15854 22330
rect 15866 22278 15918 22330
rect 15930 22278 15982 22330
rect 45122 22278 45174 22330
rect 45186 22278 45238 22330
rect 45250 22278 45302 22330
rect 45314 22278 45366 22330
rect 45378 22278 45430 22330
rect 74570 22278 74622 22330
rect 74634 22278 74686 22330
rect 74698 22278 74750 22330
rect 74762 22278 74814 22330
rect 74826 22278 74878 22330
rect 104018 22278 104070 22330
rect 104082 22278 104134 22330
rect 104146 22278 104198 22330
rect 104210 22278 104262 22330
rect 104274 22278 104326 22330
rect 50712 22083 50764 22092
rect 50712 22049 50721 22083
rect 50721 22049 50755 22083
rect 50755 22049 50764 22083
rect 50712 22040 50764 22049
rect 51080 21972 51132 22024
rect 1400 21879 1452 21888
rect 1400 21845 1409 21879
rect 1409 21845 1443 21879
rect 1443 21845 1452 21879
rect 1400 21836 1452 21845
rect 68192 21904 68244 21956
rect 50620 21879 50672 21888
rect 50620 21845 50629 21879
rect 50629 21845 50663 21879
rect 50663 21845 50672 21879
rect 50620 21836 50672 21845
rect 106372 21836 106424 21888
rect 30398 21734 30450 21786
rect 30462 21734 30514 21786
rect 30526 21734 30578 21786
rect 30590 21734 30642 21786
rect 30654 21734 30706 21786
rect 59846 21734 59898 21786
rect 59910 21734 59962 21786
rect 59974 21734 60026 21786
rect 60038 21734 60090 21786
rect 60102 21734 60154 21786
rect 89294 21734 89346 21786
rect 89358 21734 89410 21786
rect 89422 21734 89474 21786
rect 89486 21734 89538 21786
rect 89550 21734 89602 21786
rect 49700 21632 49752 21684
rect 50712 21632 50764 21684
rect 68192 21675 68244 21684
rect 68192 21641 68201 21675
rect 68201 21641 68235 21675
rect 68235 21641 68244 21675
rect 68192 21632 68244 21641
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 54484 21496 54536 21548
rect 68100 21496 68152 21548
rect 68652 21471 68704 21480
rect 68652 21437 68661 21471
rect 68661 21437 68695 21471
rect 68695 21437 68704 21471
rect 68652 21428 68704 21437
rect 68744 21471 68796 21480
rect 68744 21437 68753 21471
rect 68753 21437 68787 21471
rect 68787 21437 68796 21471
rect 68744 21428 68796 21437
rect 79232 21428 79284 21480
rect 117320 21471 117372 21480
rect 117320 21437 117329 21471
rect 117329 21437 117363 21471
rect 117363 21437 117372 21471
rect 117320 21428 117372 21437
rect 117596 21471 117648 21480
rect 117596 21437 117605 21471
rect 117605 21437 117639 21471
rect 117639 21437 117648 21471
rect 117596 21428 117648 21437
rect 28908 21360 28960 21412
rect 82728 21360 82780 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 15674 21190 15726 21242
rect 15738 21190 15790 21242
rect 15802 21190 15854 21242
rect 15866 21190 15918 21242
rect 15930 21190 15982 21242
rect 45122 21190 45174 21242
rect 45186 21190 45238 21242
rect 45250 21190 45302 21242
rect 45314 21190 45366 21242
rect 45378 21190 45430 21242
rect 74570 21190 74622 21242
rect 74634 21190 74686 21242
rect 74698 21190 74750 21242
rect 74762 21190 74814 21242
rect 74826 21190 74878 21242
rect 104018 21190 104070 21242
rect 104082 21190 104134 21242
rect 104146 21190 104198 21242
rect 104210 21190 104262 21242
rect 104274 21190 104326 21242
rect 1584 21088 1636 21140
rect 68652 21088 68704 21140
rect 55128 21020 55180 21072
rect 54576 20952 54628 21004
rect 72884 20995 72936 21004
rect 54484 20927 54536 20936
rect 54484 20893 54493 20927
rect 54493 20893 54527 20927
rect 54527 20893 54536 20927
rect 54484 20884 54536 20893
rect 55496 20884 55548 20936
rect 72884 20961 72893 20995
rect 72893 20961 72927 20995
rect 72927 20961 72936 20995
rect 72884 20952 72936 20961
rect 72700 20927 72752 20936
rect 72700 20893 72709 20927
rect 72709 20893 72743 20927
rect 72743 20893 72752 20927
rect 72700 20884 72752 20893
rect 117596 21020 117648 21072
rect 85028 20995 85080 21004
rect 85028 20961 85037 20995
rect 85037 20961 85071 20995
rect 85071 20961 85080 20995
rect 85028 20952 85080 20961
rect 115940 20884 115992 20936
rect 118056 20816 118108 20868
rect 68744 20748 68796 20800
rect 71872 20748 71924 20800
rect 72792 20791 72844 20800
rect 72792 20757 72801 20791
rect 72801 20757 72835 20791
rect 72835 20757 72844 20791
rect 84476 20791 84528 20800
rect 72792 20748 72844 20757
rect 84476 20757 84485 20791
rect 84485 20757 84519 20791
rect 84519 20757 84528 20791
rect 84476 20748 84528 20757
rect 117964 20791 118016 20800
rect 117964 20757 117973 20791
rect 117973 20757 118007 20791
rect 118007 20757 118016 20791
rect 117964 20748 118016 20757
rect 30398 20646 30450 20698
rect 30462 20646 30514 20698
rect 30526 20646 30578 20698
rect 30590 20646 30642 20698
rect 30654 20646 30706 20698
rect 59846 20646 59898 20698
rect 59910 20646 59962 20698
rect 59974 20646 60026 20698
rect 60038 20646 60090 20698
rect 60102 20646 60154 20698
rect 89294 20646 89346 20698
rect 89358 20646 89410 20698
rect 89422 20646 89474 20698
rect 89486 20646 89538 20698
rect 89550 20646 89602 20698
rect 86868 20544 86920 20596
rect 115940 20544 115992 20596
rect 71872 20451 71924 20460
rect 71872 20417 71881 20451
rect 71881 20417 71915 20451
rect 71915 20417 71924 20451
rect 71872 20408 71924 20417
rect 79048 20451 79100 20460
rect 79048 20417 79057 20451
rect 79057 20417 79091 20451
rect 79091 20417 79100 20451
rect 79048 20408 79100 20417
rect 84476 20408 84528 20460
rect 114744 20451 114796 20460
rect 114744 20417 114753 20451
rect 114753 20417 114787 20451
rect 114787 20417 114796 20451
rect 114744 20408 114796 20417
rect 79232 20383 79284 20392
rect 79232 20349 79241 20383
rect 79241 20349 79275 20383
rect 79275 20349 79284 20383
rect 79232 20340 79284 20349
rect 78036 20272 78088 20324
rect 72056 20247 72108 20256
rect 72056 20213 72065 20247
rect 72065 20213 72099 20247
rect 72099 20213 72108 20247
rect 72056 20204 72108 20213
rect 78680 20247 78732 20256
rect 78680 20213 78689 20247
rect 78689 20213 78723 20247
rect 78723 20213 78732 20247
rect 78680 20204 78732 20213
rect 15674 20102 15726 20154
rect 15738 20102 15790 20154
rect 15802 20102 15854 20154
rect 15866 20102 15918 20154
rect 15930 20102 15982 20154
rect 45122 20102 45174 20154
rect 45186 20102 45238 20154
rect 45250 20102 45302 20154
rect 45314 20102 45366 20154
rect 45378 20102 45430 20154
rect 74570 20102 74622 20154
rect 74634 20102 74686 20154
rect 74698 20102 74750 20154
rect 74762 20102 74814 20154
rect 74826 20102 74878 20154
rect 104018 20102 104070 20154
rect 104082 20102 104134 20154
rect 104146 20102 104198 20154
rect 104210 20102 104262 20154
rect 104274 20102 104326 20154
rect 47032 20000 47084 20052
rect 79048 20000 79100 20052
rect 72056 19796 72108 19848
rect 78680 19796 78732 19848
rect 78956 19728 79008 19780
rect 114744 19728 114796 19780
rect 1400 19703 1452 19712
rect 1400 19669 1409 19703
rect 1409 19669 1443 19703
rect 1443 19669 1452 19703
rect 1400 19660 1452 19669
rect 80704 19660 80756 19712
rect 113732 19703 113784 19712
rect 113732 19669 113741 19703
rect 113741 19669 113775 19703
rect 113775 19669 113784 19703
rect 113732 19660 113784 19669
rect 117964 19703 118016 19712
rect 117964 19669 117973 19703
rect 117973 19669 118007 19703
rect 118007 19669 118016 19703
rect 117964 19660 118016 19669
rect 30398 19558 30450 19610
rect 30462 19558 30514 19610
rect 30526 19558 30578 19610
rect 30590 19558 30642 19610
rect 30654 19558 30706 19610
rect 59846 19558 59898 19610
rect 59910 19558 59962 19610
rect 59974 19558 60026 19610
rect 60038 19558 60090 19610
rect 60102 19558 60154 19610
rect 89294 19558 89346 19610
rect 89358 19558 89410 19610
rect 89422 19558 89474 19610
rect 89486 19558 89538 19610
rect 89550 19558 89602 19610
rect 102692 19456 102744 19508
rect 113732 19456 113784 19508
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 66536 19116 66588 19168
rect 15674 19014 15726 19066
rect 15738 19014 15790 19066
rect 15802 19014 15854 19066
rect 15866 19014 15918 19066
rect 15930 19014 15982 19066
rect 45122 19014 45174 19066
rect 45186 19014 45238 19066
rect 45250 19014 45302 19066
rect 45314 19014 45366 19066
rect 45378 19014 45430 19066
rect 74570 19014 74622 19066
rect 74634 19014 74686 19066
rect 74698 19014 74750 19066
rect 74762 19014 74814 19066
rect 74826 19014 74878 19066
rect 104018 19014 104070 19066
rect 104082 19014 104134 19066
rect 104146 19014 104198 19066
rect 104210 19014 104262 19066
rect 104274 19014 104326 19066
rect 33324 18708 33376 18760
rect 117872 18751 117924 18760
rect 117872 18717 117881 18751
rect 117881 18717 117915 18751
rect 117915 18717 117924 18751
rect 117872 18708 117924 18717
rect 2228 18640 2280 18692
rect 68560 18640 68612 18692
rect 1400 18615 1452 18624
rect 1400 18581 1409 18615
rect 1409 18581 1443 18615
rect 1443 18581 1452 18615
rect 1400 18572 1452 18581
rect 117964 18572 118016 18624
rect 30398 18470 30450 18522
rect 30462 18470 30514 18522
rect 30526 18470 30578 18522
rect 30590 18470 30642 18522
rect 30654 18470 30706 18522
rect 59846 18470 59898 18522
rect 59910 18470 59962 18522
rect 59974 18470 60026 18522
rect 60038 18470 60090 18522
rect 60102 18470 60154 18522
rect 89294 18470 89346 18522
rect 89358 18470 89410 18522
rect 89422 18470 89474 18522
rect 89486 18470 89538 18522
rect 89550 18470 89602 18522
rect 33324 18275 33376 18284
rect 33324 18241 33333 18275
rect 33333 18241 33367 18275
rect 33367 18241 33376 18275
rect 33324 18232 33376 18241
rect 117872 18275 117924 18284
rect 117872 18241 117881 18275
rect 117881 18241 117915 18275
rect 117915 18241 117924 18275
rect 117872 18232 117924 18241
rect 33232 18164 33284 18216
rect 117688 18028 117740 18080
rect 15674 17926 15726 17978
rect 15738 17926 15790 17978
rect 15802 17926 15854 17978
rect 15866 17926 15918 17978
rect 15930 17926 15982 17978
rect 45122 17926 45174 17978
rect 45186 17926 45238 17978
rect 45250 17926 45302 17978
rect 45314 17926 45366 17978
rect 45378 17926 45430 17978
rect 74570 17926 74622 17978
rect 74634 17926 74686 17978
rect 74698 17926 74750 17978
rect 74762 17926 74814 17978
rect 74826 17926 74878 17978
rect 104018 17926 104070 17978
rect 104082 17926 104134 17978
rect 104146 17926 104198 17978
rect 104210 17926 104262 17978
rect 104274 17926 104326 17978
rect 33232 17824 33284 17876
rect 81440 17756 81492 17808
rect 82728 17756 82780 17808
rect 31300 17688 31352 17740
rect 37832 17688 37884 17740
rect 26884 17620 26936 17672
rect 33784 17527 33836 17536
rect 33784 17493 33793 17527
rect 33793 17493 33827 17527
rect 33827 17493 33836 17527
rect 33784 17484 33836 17493
rect 30398 17382 30450 17434
rect 30462 17382 30514 17434
rect 30526 17382 30578 17434
rect 30590 17382 30642 17434
rect 30654 17382 30706 17434
rect 59846 17382 59898 17434
rect 59910 17382 59962 17434
rect 59974 17382 60026 17434
rect 60038 17382 60090 17434
rect 60102 17382 60154 17434
rect 89294 17382 89346 17434
rect 89358 17382 89410 17434
rect 89422 17382 89474 17434
rect 89486 17382 89538 17434
rect 89550 17382 89602 17434
rect 59728 17280 59780 17332
rect 70124 17280 70176 17332
rect 65984 17212 66036 17264
rect 115204 17212 115256 17264
rect 1952 17144 2004 17196
rect 82912 17187 82964 17196
rect 82912 17153 82921 17187
rect 82921 17153 82955 17187
rect 82955 17153 82964 17187
rect 82912 17144 82964 17153
rect 1400 17051 1452 17060
rect 1400 17017 1409 17051
rect 1409 17017 1443 17051
rect 1443 17017 1452 17051
rect 1400 17008 1452 17017
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 90364 16940 90416 16992
rect 15674 16838 15726 16890
rect 15738 16838 15790 16890
rect 15802 16838 15854 16890
rect 15866 16838 15918 16890
rect 15930 16838 15982 16890
rect 45122 16838 45174 16890
rect 45186 16838 45238 16890
rect 45250 16838 45302 16890
rect 45314 16838 45366 16890
rect 45378 16838 45430 16890
rect 74570 16838 74622 16890
rect 74634 16838 74686 16890
rect 74698 16838 74750 16890
rect 74762 16838 74814 16890
rect 74826 16838 74878 16890
rect 104018 16838 104070 16890
rect 104082 16838 104134 16890
rect 104146 16838 104198 16890
rect 104210 16838 104262 16890
rect 104274 16838 104326 16890
rect 25412 16668 25464 16720
rect 3516 16600 3568 16652
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 70584 16532 70636 16584
rect 82728 16643 82780 16652
rect 82728 16609 82737 16643
rect 82737 16609 82771 16643
rect 82771 16609 82780 16643
rect 82728 16600 82780 16609
rect 2596 16464 2648 16516
rect 70768 16464 70820 16516
rect 117228 16532 117280 16584
rect 1952 16396 2004 16448
rect 82912 16396 82964 16448
rect 30398 16294 30450 16346
rect 30462 16294 30514 16346
rect 30526 16294 30578 16346
rect 30590 16294 30642 16346
rect 30654 16294 30706 16346
rect 59846 16294 59898 16346
rect 59910 16294 59962 16346
rect 59974 16294 60026 16346
rect 60038 16294 60090 16346
rect 60102 16294 60154 16346
rect 89294 16294 89346 16346
rect 89358 16294 89410 16346
rect 89422 16294 89474 16346
rect 89486 16294 89538 16346
rect 89550 16294 89602 16346
rect 68284 16124 68336 16176
rect 67456 16056 67508 16108
rect 68468 16056 68520 16108
rect 69572 16056 69624 16108
rect 68928 15920 68980 15972
rect 68376 15852 68428 15904
rect 70584 15852 70636 15904
rect 118148 15895 118200 15904
rect 118148 15861 118157 15895
rect 118157 15861 118191 15895
rect 118191 15861 118200 15895
rect 118148 15852 118200 15861
rect 15674 15750 15726 15802
rect 15738 15750 15790 15802
rect 15802 15750 15854 15802
rect 15866 15750 15918 15802
rect 15930 15750 15982 15802
rect 45122 15750 45174 15802
rect 45186 15750 45238 15802
rect 45250 15750 45302 15802
rect 45314 15750 45366 15802
rect 45378 15750 45430 15802
rect 74570 15750 74622 15802
rect 74634 15750 74686 15802
rect 74698 15750 74750 15802
rect 74762 15750 74814 15802
rect 74826 15750 74878 15802
rect 104018 15750 104070 15802
rect 104082 15750 104134 15802
rect 104146 15750 104198 15802
rect 104210 15750 104262 15802
rect 104274 15750 104326 15802
rect 53840 15512 53892 15564
rect 67088 15512 67140 15564
rect 68836 15648 68888 15700
rect 69572 15691 69624 15700
rect 69572 15657 69581 15691
rect 69581 15657 69615 15691
rect 69615 15657 69624 15691
rect 69572 15648 69624 15657
rect 70768 15691 70820 15700
rect 70768 15657 70777 15691
rect 70777 15657 70811 15691
rect 70811 15657 70820 15691
rect 70768 15648 70820 15657
rect 68284 15555 68336 15564
rect 68284 15521 68293 15555
rect 68293 15521 68327 15555
rect 68327 15521 68336 15555
rect 71320 15555 71372 15564
rect 68284 15512 68336 15521
rect 71320 15521 71329 15555
rect 71329 15521 71363 15555
rect 71363 15521 71372 15555
rect 71320 15512 71372 15521
rect 10416 15444 10468 15496
rect 1400 15351 1452 15360
rect 1400 15317 1409 15351
rect 1409 15317 1443 15351
rect 1443 15317 1452 15351
rect 1400 15308 1452 15317
rect 10876 15308 10928 15360
rect 56692 15444 56744 15496
rect 64972 15444 65024 15496
rect 65984 15487 66036 15496
rect 65984 15453 65993 15487
rect 65993 15453 66027 15487
rect 66027 15453 66036 15487
rect 65984 15444 66036 15453
rect 67180 15487 67232 15496
rect 67180 15453 67189 15487
rect 67189 15453 67223 15487
rect 67223 15453 67232 15487
rect 67180 15444 67232 15453
rect 67732 15444 67784 15496
rect 68192 15487 68244 15496
rect 68192 15453 68201 15487
rect 68201 15453 68235 15487
rect 68235 15453 68244 15487
rect 68192 15444 68244 15453
rect 69204 15487 69256 15496
rect 32772 15308 32824 15360
rect 64696 15351 64748 15360
rect 64696 15317 64705 15351
rect 64705 15317 64739 15351
rect 64739 15317 64748 15351
rect 64696 15308 64748 15317
rect 65800 15308 65852 15360
rect 66996 15351 67048 15360
rect 66996 15317 67005 15351
rect 67005 15317 67039 15351
rect 67039 15317 67048 15351
rect 66996 15308 67048 15317
rect 67548 15308 67600 15360
rect 69204 15453 69213 15487
rect 69213 15453 69247 15487
rect 69247 15453 69256 15487
rect 69204 15444 69256 15453
rect 68744 15376 68796 15428
rect 69664 15376 69716 15428
rect 117412 15376 117464 15428
rect 69756 15308 69808 15360
rect 71136 15351 71188 15360
rect 71136 15317 71145 15351
rect 71145 15317 71179 15351
rect 71179 15317 71188 15351
rect 71136 15308 71188 15317
rect 112536 15308 112588 15360
rect 30398 15206 30450 15258
rect 30462 15206 30514 15258
rect 30526 15206 30578 15258
rect 30590 15206 30642 15258
rect 30654 15206 30706 15258
rect 59846 15206 59898 15258
rect 59910 15206 59962 15258
rect 59974 15206 60026 15258
rect 60038 15206 60090 15258
rect 60102 15206 60154 15258
rect 89294 15206 89346 15258
rect 89358 15206 89410 15258
rect 89422 15206 89474 15258
rect 89486 15206 89538 15258
rect 89550 15206 89602 15258
rect 10416 15104 10468 15156
rect 64880 15104 64932 15156
rect 118056 15104 118108 15156
rect 64144 15036 64196 15088
rect 65064 15036 65116 15088
rect 66536 15079 66588 15088
rect 66536 15045 66545 15079
rect 66545 15045 66579 15079
rect 66579 15045 66588 15079
rect 66536 15036 66588 15045
rect 68744 15079 68796 15088
rect 68744 15045 68753 15079
rect 68753 15045 68787 15079
rect 68787 15045 68796 15079
rect 68744 15036 68796 15045
rect 68836 15036 68888 15088
rect 69664 15036 69716 15088
rect 70584 15036 70636 15088
rect 2412 14968 2464 15020
rect 10876 14968 10928 15020
rect 50528 14968 50580 15020
rect 64696 14968 64748 15020
rect 65892 15011 65944 15020
rect 65892 14977 65901 15011
rect 65901 14977 65935 15011
rect 65935 14977 65944 15011
rect 65892 14968 65944 14977
rect 69204 15011 69256 15020
rect 41328 14900 41380 14952
rect 54576 14943 54628 14952
rect 54576 14909 54585 14943
rect 54585 14909 54619 14943
rect 54619 14909 54628 14943
rect 54576 14900 54628 14909
rect 56140 14943 56192 14952
rect 56140 14909 56149 14943
rect 56149 14909 56183 14943
rect 56183 14909 56192 14943
rect 56140 14900 56192 14909
rect 64144 14900 64196 14952
rect 43352 14832 43404 14884
rect 64972 14832 65024 14884
rect 68468 14900 68520 14952
rect 68652 14832 68704 14884
rect 68836 14832 68888 14884
rect 69204 14977 69213 15011
rect 69213 14977 69247 15011
rect 69247 14977 69256 15011
rect 69204 14968 69256 14977
rect 69296 15011 69348 15020
rect 69296 14977 69305 15011
rect 69305 14977 69339 15011
rect 69339 14977 69348 15011
rect 69296 14968 69348 14977
rect 70400 14968 70452 15020
rect 71228 15036 71280 15088
rect 70032 14943 70084 14952
rect 70032 14909 70041 14943
rect 70041 14909 70075 14943
rect 70075 14909 70084 14943
rect 70032 14900 70084 14909
rect 69296 14832 69348 14884
rect 37832 14764 37884 14816
rect 53840 14807 53892 14816
rect 53840 14773 53849 14807
rect 53849 14773 53883 14807
rect 53883 14773 53892 14807
rect 53840 14764 53892 14773
rect 58532 14764 58584 14816
rect 65984 14807 66036 14816
rect 65984 14773 65993 14807
rect 65993 14773 66027 14807
rect 66027 14773 66036 14807
rect 65984 14764 66036 14773
rect 66076 14764 66128 14816
rect 69020 14764 69072 14816
rect 69848 14764 69900 14816
rect 70216 14832 70268 14884
rect 94964 14900 95016 14952
rect 70308 14807 70360 14816
rect 70308 14773 70317 14807
rect 70317 14773 70351 14807
rect 70351 14773 70360 14807
rect 70308 14764 70360 14773
rect 70584 14764 70636 14816
rect 15674 14662 15726 14714
rect 15738 14662 15790 14714
rect 15802 14662 15854 14714
rect 15866 14662 15918 14714
rect 15930 14662 15982 14714
rect 45122 14662 45174 14714
rect 45186 14662 45238 14714
rect 45250 14662 45302 14714
rect 45314 14662 45366 14714
rect 45378 14662 45430 14714
rect 74570 14662 74622 14714
rect 74634 14662 74686 14714
rect 74698 14662 74750 14714
rect 74762 14662 74814 14714
rect 74826 14662 74878 14714
rect 104018 14662 104070 14714
rect 104082 14662 104134 14714
rect 104146 14662 104198 14714
rect 104210 14662 104262 14714
rect 104274 14662 104326 14714
rect 55496 14603 55548 14612
rect 55496 14569 55505 14603
rect 55505 14569 55539 14603
rect 55539 14569 55548 14603
rect 55496 14560 55548 14569
rect 67088 14560 67140 14612
rect 118056 14603 118108 14612
rect 118056 14569 118065 14603
rect 118065 14569 118099 14603
rect 118099 14569 118108 14603
rect 118056 14560 118108 14569
rect 69848 14492 69900 14544
rect 71412 14492 71464 14544
rect 50436 14424 50488 14476
rect 2412 14399 2464 14408
rect 2412 14365 2421 14399
rect 2421 14365 2455 14399
rect 2455 14365 2464 14399
rect 2412 14356 2464 14365
rect 50528 14356 50580 14408
rect 54576 14356 54628 14408
rect 1400 14263 1452 14272
rect 1400 14229 1409 14263
rect 1409 14229 1443 14263
rect 1443 14229 1452 14263
rect 1400 14220 1452 14229
rect 50804 14220 50856 14272
rect 65892 14356 65944 14408
rect 66076 14288 66128 14340
rect 64972 14220 65024 14272
rect 69664 14424 69716 14476
rect 68652 14399 68704 14408
rect 68652 14365 68661 14399
rect 68661 14365 68695 14399
rect 68695 14365 68704 14399
rect 68652 14356 68704 14365
rect 71044 14399 71096 14408
rect 67824 14288 67876 14340
rect 68928 14331 68980 14340
rect 68928 14297 68962 14331
rect 68962 14297 68980 14331
rect 68928 14288 68980 14297
rect 69020 14288 69072 14340
rect 70584 14288 70636 14340
rect 70676 14288 70728 14340
rect 71044 14365 71053 14399
rect 71053 14365 71087 14399
rect 71087 14365 71096 14399
rect 71044 14356 71096 14365
rect 71504 14399 71556 14408
rect 71504 14365 71513 14399
rect 71513 14365 71547 14399
rect 71547 14365 71556 14399
rect 71504 14356 71556 14365
rect 117872 14399 117924 14408
rect 117872 14365 117881 14399
rect 117881 14365 117915 14399
rect 117915 14365 117924 14399
rect 117872 14356 117924 14365
rect 90640 14288 90692 14340
rect 68468 14220 68520 14272
rect 69296 14220 69348 14272
rect 70400 14220 70452 14272
rect 30398 14118 30450 14170
rect 30462 14118 30514 14170
rect 30526 14118 30578 14170
rect 30590 14118 30642 14170
rect 30654 14118 30706 14170
rect 59846 14118 59898 14170
rect 59910 14118 59962 14170
rect 59974 14118 60026 14170
rect 60038 14118 60090 14170
rect 60102 14118 60154 14170
rect 89294 14118 89346 14170
rect 89358 14118 89410 14170
rect 89422 14118 89474 14170
rect 89486 14118 89538 14170
rect 89550 14118 89602 14170
rect 56140 14016 56192 14068
rect 65984 14016 66036 14068
rect 67180 14016 67232 14068
rect 69020 14016 69072 14068
rect 65800 13923 65852 13932
rect 65800 13889 65809 13923
rect 65809 13889 65843 13923
rect 65843 13889 65852 13923
rect 65800 13880 65852 13889
rect 69664 13948 69716 14000
rect 69756 13948 69808 14000
rect 71412 14016 71464 14068
rect 86224 14059 86276 14068
rect 86224 14025 86233 14059
rect 86233 14025 86267 14059
rect 86267 14025 86276 14059
rect 86224 14016 86276 14025
rect 118240 14016 118292 14068
rect 86408 13948 86460 14000
rect 68560 13923 68612 13932
rect 66260 13855 66312 13864
rect 66260 13821 66269 13855
rect 66269 13821 66303 13855
rect 66303 13821 66312 13855
rect 66260 13812 66312 13821
rect 68560 13889 68569 13923
rect 68569 13889 68603 13923
rect 68603 13889 68612 13923
rect 68560 13880 68612 13889
rect 68836 13880 68888 13932
rect 70676 13880 70728 13932
rect 71504 13880 71556 13932
rect 69572 13812 69624 13864
rect 69848 13812 69900 13864
rect 70768 13855 70820 13864
rect 70768 13821 70777 13855
rect 70777 13821 70811 13855
rect 70811 13821 70820 13855
rect 70768 13812 70820 13821
rect 81992 13812 82044 13864
rect 86316 13855 86368 13864
rect 86316 13821 86325 13855
rect 86325 13821 86359 13855
rect 86359 13821 86368 13855
rect 86316 13812 86368 13821
rect 86408 13855 86460 13864
rect 86408 13821 86417 13855
rect 86417 13821 86451 13855
rect 86451 13821 86460 13855
rect 108120 13880 108172 13932
rect 117872 13923 117924 13932
rect 117872 13889 117881 13923
rect 117881 13889 117915 13923
rect 117915 13889 117924 13923
rect 117872 13880 117924 13889
rect 86408 13812 86460 13821
rect 48504 13744 48556 13796
rect 57612 13744 57664 13796
rect 70400 13744 70452 13796
rect 68192 13676 68244 13728
rect 68744 13676 68796 13728
rect 69848 13719 69900 13728
rect 69848 13685 69857 13719
rect 69857 13685 69891 13719
rect 69891 13685 69900 13719
rect 69848 13676 69900 13685
rect 86776 13676 86828 13728
rect 15674 13574 15726 13626
rect 15738 13574 15790 13626
rect 15802 13574 15854 13626
rect 15866 13574 15918 13626
rect 15930 13574 15982 13626
rect 45122 13574 45174 13626
rect 45186 13574 45238 13626
rect 45250 13574 45302 13626
rect 45314 13574 45366 13626
rect 45378 13574 45430 13626
rect 74570 13574 74622 13626
rect 74634 13574 74686 13626
rect 74698 13574 74750 13626
rect 74762 13574 74814 13626
rect 74826 13574 74878 13626
rect 104018 13574 104070 13626
rect 104082 13574 104134 13626
rect 104146 13574 104198 13626
rect 104210 13574 104262 13626
rect 104274 13574 104326 13626
rect 68652 13472 68704 13524
rect 70032 13472 70084 13524
rect 69020 13268 69072 13320
rect 69848 13268 69900 13320
rect 86776 13311 86828 13320
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 16028 13200 16080 13252
rect 42984 13200 43036 13252
rect 67732 13200 67784 13252
rect 86776 13277 86785 13311
rect 86785 13277 86819 13311
rect 86819 13277 86828 13311
rect 86776 13268 86828 13277
rect 118148 13311 118200 13320
rect 118148 13277 118157 13311
rect 118157 13277 118191 13311
rect 118191 13277 118200 13311
rect 118148 13268 118200 13277
rect 31116 13132 31168 13184
rect 86592 13175 86644 13184
rect 86592 13141 86601 13175
rect 86601 13141 86635 13175
rect 86635 13141 86644 13175
rect 86592 13132 86644 13141
rect 117964 13175 118016 13184
rect 117964 13141 117973 13175
rect 117973 13141 118007 13175
rect 118007 13141 118016 13175
rect 117964 13132 118016 13141
rect 30398 13030 30450 13082
rect 30462 13030 30514 13082
rect 30526 13030 30578 13082
rect 30590 13030 30642 13082
rect 30654 13030 30706 13082
rect 59846 13030 59898 13082
rect 59910 13030 59962 13082
rect 59974 13030 60026 13082
rect 60038 13030 60090 13082
rect 60102 13030 60154 13082
rect 89294 13030 89346 13082
rect 89358 13030 89410 13082
rect 89422 13030 89474 13082
rect 89486 13030 89538 13082
rect 89550 13030 89602 13082
rect 32128 12971 32180 12980
rect 32128 12937 32137 12971
rect 32137 12937 32171 12971
rect 32171 12937 32180 12971
rect 32128 12928 32180 12937
rect 67732 12928 67784 12980
rect 67824 12928 67876 12980
rect 71044 12928 71096 12980
rect 73804 12928 73856 12980
rect 66996 12860 67048 12912
rect 20628 12792 20680 12844
rect 32312 12835 32364 12844
rect 32312 12801 32321 12835
rect 32321 12801 32355 12835
rect 32355 12801 32364 12835
rect 32312 12792 32364 12801
rect 66260 12835 66312 12844
rect 66260 12801 66269 12835
rect 66269 12801 66303 12835
rect 66303 12801 66312 12835
rect 66260 12792 66312 12801
rect 68376 12835 68428 12844
rect 68376 12801 68385 12835
rect 68385 12801 68419 12835
rect 68419 12801 68428 12835
rect 68376 12792 68428 12801
rect 70308 12860 70360 12912
rect 68744 12792 68796 12844
rect 108120 12792 108172 12844
rect 67272 12724 67324 12776
rect 68836 12724 68888 12776
rect 77024 12767 77076 12776
rect 77024 12733 77033 12767
rect 77033 12733 77067 12767
rect 77067 12733 77076 12767
rect 77024 12724 77076 12733
rect 1400 12631 1452 12640
rect 1400 12597 1409 12631
rect 1409 12597 1443 12631
rect 1443 12597 1452 12631
rect 1400 12588 1452 12597
rect 68284 12588 68336 12640
rect 76380 12631 76432 12640
rect 76380 12597 76389 12631
rect 76389 12597 76423 12631
rect 76423 12597 76432 12631
rect 76380 12588 76432 12597
rect 99380 12588 99432 12640
rect 118148 12588 118200 12640
rect 15674 12486 15726 12538
rect 15738 12486 15790 12538
rect 15802 12486 15854 12538
rect 15866 12486 15918 12538
rect 15930 12486 15982 12538
rect 45122 12486 45174 12538
rect 45186 12486 45238 12538
rect 45250 12486 45302 12538
rect 45314 12486 45366 12538
rect 45378 12486 45430 12538
rect 74570 12486 74622 12538
rect 74634 12486 74686 12538
rect 74698 12486 74750 12538
rect 74762 12486 74814 12538
rect 74826 12486 74878 12538
rect 104018 12486 104070 12538
rect 104082 12486 104134 12538
rect 104146 12486 104198 12538
rect 104210 12486 104262 12538
rect 104274 12486 104326 12538
rect 20628 12384 20680 12436
rect 32312 12384 32364 12436
rect 67180 12384 67232 12436
rect 67456 12427 67508 12436
rect 67456 12393 67465 12427
rect 67465 12393 67499 12427
rect 67499 12393 67508 12427
rect 67456 12384 67508 12393
rect 68284 12427 68336 12436
rect 68284 12393 68293 12427
rect 68293 12393 68327 12427
rect 68327 12393 68336 12427
rect 68284 12384 68336 12393
rect 11704 12248 11756 12300
rect 39396 12316 39448 12368
rect 41328 12316 41380 12368
rect 29736 12180 29788 12232
rect 55496 12180 55548 12232
rect 70768 12180 70820 12232
rect 71688 12180 71740 12232
rect 23296 12112 23348 12164
rect 43996 12155 44048 12164
rect 43996 12121 44005 12155
rect 44005 12121 44039 12155
rect 44039 12121 44048 12155
rect 43996 12112 44048 12121
rect 67088 12155 67140 12164
rect 67088 12121 67097 12155
rect 67097 12121 67131 12155
rect 67131 12121 67140 12155
rect 67088 12112 67140 12121
rect 67548 12112 67600 12164
rect 30840 12087 30892 12096
rect 30840 12053 30849 12087
rect 30849 12053 30883 12087
rect 30883 12053 30892 12087
rect 30840 12044 30892 12053
rect 71412 12044 71464 12096
rect 87236 12044 87288 12096
rect 30398 11942 30450 11994
rect 30462 11942 30514 11994
rect 30526 11942 30578 11994
rect 30590 11942 30642 11994
rect 30654 11942 30706 11994
rect 59846 11942 59898 11994
rect 59910 11942 59962 11994
rect 59974 11942 60026 11994
rect 60038 11942 60090 11994
rect 60102 11942 60154 11994
rect 89294 11942 89346 11994
rect 89358 11942 89410 11994
rect 89422 11942 89474 11994
rect 89486 11942 89538 11994
rect 89550 11942 89602 11994
rect 7840 11840 7892 11892
rect 30840 11840 30892 11892
rect 38476 11840 38528 11892
rect 75552 11840 75604 11892
rect 95240 11840 95292 11892
rect 76380 11772 76432 11824
rect 1492 11704 1544 11756
rect 71688 11704 71740 11756
rect 99656 11772 99708 11824
rect 1400 11611 1452 11620
rect 1400 11577 1409 11611
rect 1409 11577 1443 11611
rect 1443 11577 1452 11611
rect 1400 11568 1452 11577
rect 39396 11679 39448 11688
rect 39396 11645 39405 11679
rect 39405 11645 39439 11679
rect 39439 11645 39448 11679
rect 39396 11636 39448 11645
rect 43996 11636 44048 11688
rect 77024 11636 77076 11688
rect 117320 11679 117372 11688
rect 117320 11645 117329 11679
rect 117329 11645 117363 11679
rect 117363 11645 117372 11679
rect 117320 11636 117372 11645
rect 117412 11636 117464 11688
rect 38476 11543 38528 11552
rect 38476 11509 38485 11543
rect 38485 11509 38519 11543
rect 38519 11509 38528 11543
rect 38476 11500 38528 11509
rect 42524 11500 42576 11552
rect 118148 11500 118200 11552
rect 15674 11398 15726 11450
rect 15738 11398 15790 11450
rect 15802 11398 15854 11450
rect 15866 11398 15918 11450
rect 15930 11398 15982 11450
rect 45122 11398 45174 11450
rect 45186 11398 45238 11450
rect 45250 11398 45302 11450
rect 45314 11398 45366 11450
rect 45378 11398 45430 11450
rect 74570 11398 74622 11450
rect 74634 11398 74686 11450
rect 74698 11398 74750 11450
rect 74762 11398 74814 11450
rect 74826 11398 74878 11450
rect 104018 11398 104070 11450
rect 104082 11398 104134 11450
rect 104146 11398 104198 11450
rect 104210 11398 104262 11450
rect 104274 11398 104326 11450
rect 117964 11271 118016 11280
rect 117964 11237 117973 11271
rect 117973 11237 118007 11271
rect 118007 11237 118016 11271
rect 117964 11228 118016 11237
rect 9220 11203 9272 11212
rect 9220 11169 9229 11203
rect 9229 11169 9263 11203
rect 9263 11169 9272 11203
rect 9220 11160 9272 11169
rect 42524 11203 42576 11212
rect 42524 11169 42533 11203
rect 42533 11169 42567 11203
rect 42567 11169 42576 11203
rect 42524 11160 42576 11169
rect 2688 11092 2740 11144
rect 63408 11092 63460 11144
rect 118148 11135 118200 11144
rect 118148 11101 118157 11135
rect 118157 11101 118191 11135
rect 118191 11101 118200 11135
rect 118148 11092 118200 11101
rect 30398 10854 30450 10906
rect 30462 10854 30514 10906
rect 30526 10854 30578 10906
rect 30590 10854 30642 10906
rect 30654 10854 30706 10906
rect 59846 10854 59898 10906
rect 59910 10854 59962 10906
rect 59974 10854 60026 10906
rect 60038 10854 60090 10906
rect 60102 10854 60154 10906
rect 89294 10854 89346 10906
rect 89358 10854 89410 10906
rect 89422 10854 89474 10906
rect 89486 10854 89538 10906
rect 89550 10854 89602 10906
rect 66260 10752 66312 10804
rect 30932 10684 30984 10736
rect 2504 10616 2556 10668
rect 69020 10684 69072 10736
rect 82544 10684 82596 10736
rect 36544 10548 36596 10600
rect 91928 10548 91980 10600
rect 32956 10480 33008 10532
rect 105544 10480 105596 10532
rect 1400 10455 1452 10464
rect 1400 10421 1409 10455
rect 1409 10421 1443 10455
rect 1443 10421 1452 10455
rect 1400 10412 1452 10421
rect 83004 10412 83056 10464
rect 111708 10412 111760 10464
rect 15674 10310 15726 10362
rect 15738 10310 15790 10362
rect 15802 10310 15854 10362
rect 15866 10310 15918 10362
rect 15930 10310 15982 10362
rect 45122 10310 45174 10362
rect 45186 10310 45238 10362
rect 45250 10310 45302 10362
rect 45314 10310 45366 10362
rect 45378 10310 45430 10362
rect 74570 10310 74622 10362
rect 74634 10310 74686 10362
rect 74698 10310 74750 10362
rect 74762 10310 74814 10362
rect 74826 10310 74878 10362
rect 104018 10310 104070 10362
rect 104082 10310 104134 10362
rect 104146 10310 104198 10362
rect 104210 10310 104262 10362
rect 104274 10310 104326 10362
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 113640 10208 113692 10260
rect 1492 10004 1544 10056
rect 2688 10047 2740 10056
rect 2688 10013 2697 10047
rect 2697 10013 2731 10047
rect 2731 10013 2740 10047
rect 2688 10004 2740 10013
rect 115940 10004 115992 10056
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 1860 9936 1912 9945
rect 114744 9936 114796 9988
rect 31760 9868 31812 9920
rect 117964 9911 118016 9920
rect 117964 9877 117973 9911
rect 117973 9877 118007 9911
rect 118007 9877 118016 9911
rect 117964 9868 118016 9877
rect 30398 9766 30450 9818
rect 30462 9766 30514 9818
rect 30526 9766 30578 9818
rect 30590 9766 30642 9818
rect 30654 9766 30706 9818
rect 59846 9766 59898 9818
rect 59910 9766 59962 9818
rect 59974 9766 60026 9818
rect 60038 9766 60090 9818
rect 60102 9766 60154 9818
rect 89294 9766 89346 9818
rect 89358 9766 89410 9818
rect 89422 9766 89474 9818
rect 89486 9766 89538 9818
rect 89550 9766 89602 9818
rect 68560 9596 68612 9648
rect 115388 9596 115440 9648
rect 114744 9571 114796 9580
rect 114744 9537 114753 9571
rect 114753 9537 114787 9571
rect 114787 9537 114796 9571
rect 114744 9528 114796 9537
rect 115940 9392 115992 9444
rect 15674 9222 15726 9274
rect 15738 9222 15790 9274
rect 15802 9222 15854 9274
rect 15866 9222 15918 9274
rect 15930 9222 15982 9274
rect 45122 9222 45174 9274
rect 45186 9222 45238 9274
rect 45250 9222 45302 9274
rect 45314 9222 45366 9274
rect 45378 9222 45430 9274
rect 74570 9222 74622 9274
rect 74634 9222 74686 9274
rect 74698 9222 74750 9274
rect 74762 9222 74814 9274
rect 74826 9222 74878 9274
rect 104018 9222 104070 9274
rect 104082 9222 104134 9274
rect 104146 9222 104198 9274
rect 104210 9222 104262 9274
rect 104274 9222 104326 9274
rect 76656 8916 76708 8968
rect 113640 8916 113692 8968
rect 30398 8678 30450 8730
rect 30462 8678 30514 8730
rect 30526 8678 30578 8730
rect 30590 8678 30642 8730
rect 30654 8678 30706 8730
rect 59846 8678 59898 8730
rect 59910 8678 59962 8730
rect 59974 8678 60026 8730
rect 60038 8678 60090 8730
rect 60102 8678 60154 8730
rect 89294 8678 89346 8730
rect 89358 8678 89410 8730
rect 89422 8678 89474 8730
rect 89486 8678 89538 8730
rect 89550 8678 89602 8730
rect 77208 8440 77260 8492
rect 29460 8415 29512 8424
rect 29460 8381 29469 8415
rect 29469 8381 29503 8415
rect 29503 8381 29512 8415
rect 29460 8372 29512 8381
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 117964 8347 118016 8356
rect 117964 8313 117973 8347
rect 117973 8313 118007 8347
rect 118007 8313 118016 8347
rect 117964 8304 118016 8313
rect 15674 8134 15726 8186
rect 15738 8134 15790 8186
rect 15802 8134 15854 8186
rect 15866 8134 15918 8186
rect 15930 8134 15982 8186
rect 45122 8134 45174 8186
rect 45186 8134 45238 8186
rect 45250 8134 45302 8186
rect 45314 8134 45366 8186
rect 45378 8134 45430 8186
rect 74570 8134 74622 8186
rect 74634 8134 74686 8186
rect 74698 8134 74750 8186
rect 74762 8134 74814 8186
rect 74826 8134 74878 8186
rect 104018 8134 104070 8186
rect 104082 8134 104134 8186
rect 104146 8134 104198 8186
rect 104210 8134 104262 8186
rect 104274 8134 104326 8186
rect 29460 8032 29512 8084
rect 77208 8007 77260 8016
rect 77208 7973 77217 8007
rect 77217 7973 77251 8007
rect 77251 7973 77260 8007
rect 77208 7964 77260 7973
rect 27528 7896 27580 7948
rect 43996 7896 44048 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 46940 7760 46992 7812
rect 76472 7760 76524 7812
rect 116216 7760 116268 7812
rect 48320 7692 48372 7744
rect 30398 7590 30450 7642
rect 30462 7590 30514 7642
rect 30526 7590 30578 7642
rect 30590 7590 30642 7642
rect 30654 7590 30706 7642
rect 59846 7590 59898 7642
rect 59910 7590 59962 7642
rect 59974 7590 60026 7642
rect 60038 7590 60090 7642
rect 60102 7590 60154 7642
rect 89294 7590 89346 7642
rect 89358 7590 89410 7642
rect 89422 7590 89474 7642
rect 89486 7590 89538 7642
rect 89550 7590 89602 7642
rect 70492 7488 70544 7540
rect 71320 7488 71372 7540
rect 86960 7352 87012 7404
rect 117964 7395 118016 7404
rect 117964 7361 117973 7395
rect 117973 7361 118007 7395
rect 118007 7361 118016 7395
rect 117964 7352 118016 7361
rect 4804 7148 4856 7200
rect 86960 7148 87012 7200
rect 15674 7046 15726 7098
rect 15738 7046 15790 7098
rect 15802 7046 15854 7098
rect 15866 7046 15918 7098
rect 15930 7046 15982 7098
rect 45122 7046 45174 7098
rect 45186 7046 45238 7098
rect 45250 7046 45302 7098
rect 45314 7046 45366 7098
rect 45378 7046 45430 7098
rect 74570 7046 74622 7098
rect 74634 7046 74686 7098
rect 74698 7046 74750 7098
rect 74762 7046 74814 7098
rect 74826 7046 74878 7098
rect 104018 7046 104070 7098
rect 104082 7046 104134 7098
rect 104146 7046 104198 7098
rect 104210 7046 104262 7098
rect 104274 7046 104326 7098
rect 64604 6876 64656 6928
rect 69480 6876 69532 6928
rect 49884 6740 49936 6792
rect 50068 6604 50120 6656
rect 30398 6502 30450 6554
rect 30462 6502 30514 6554
rect 30526 6502 30578 6554
rect 30590 6502 30642 6554
rect 30654 6502 30706 6554
rect 59846 6502 59898 6554
rect 59910 6502 59962 6554
rect 59974 6502 60026 6554
rect 60038 6502 60090 6554
rect 60102 6502 60154 6554
rect 89294 6502 89346 6554
rect 89358 6502 89410 6554
rect 89422 6502 89474 6554
rect 89486 6502 89538 6554
rect 89550 6502 89602 6554
rect 49884 6443 49936 6452
rect 49884 6409 49893 6443
rect 49893 6409 49927 6443
rect 49927 6409 49936 6443
rect 49884 6400 49936 6409
rect 1952 6264 2004 6316
rect 49700 6264 49752 6316
rect 86960 6307 87012 6316
rect 50436 6239 50488 6248
rect 50436 6205 50445 6239
rect 50445 6205 50479 6239
rect 50479 6205 50488 6239
rect 86960 6273 86969 6307
rect 86969 6273 87003 6307
rect 87003 6273 87012 6307
rect 86960 6264 87012 6273
rect 117872 6307 117924 6316
rect 117872 6273 117881 6307
rect 117881 6273 117915 6307
rect 117915 6273 117924 6307
rect 117872 6264 117924 6273
rect 50436 6196 50488 6205
rect 1400 6171 1452 6180
rect 1400 6137 1409 6171
rect 1409 6137 1443 6171
rect 1443 6137 1452 6171
rect 1400 6128 1452 6137
rect 59268 6128 59320 6180
rect 110052 6128 110104 6180
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 87236 6060 87288 6112
rect 15674 5958 15726 6010
rect 15738 5958 15790 6010
rect 15802 5958 15854 6010
rect 15866 5958 15918 6010
rect 15930 5958 15982 6010
rect 45122 5958 45174 6010
rect 45186 5958 45238 6010
rect 45250 5958 45302 6010
rect 45314 5958 45366 6010
rect 45378 5958 45430 6010
rect 74570 5958 74622 6010
rect 74634 5958 74686 6010
rect 74698 5958 74750 6010
rect 74762 5958 74814 6010
rect 74826 5958 74878 6010
rect 104018 5958 104070 6010
rect 104082 5958 104134 6010
rect 104146 5958 104198 6010
rect 104210 5958 104262 6010
rect 104274 5958 104326 6010
rect 57428 5652 57480 5704
rect 65892 5652 65944 5704
rect 1860 5627 1912 5636
rect 1860 5593 1869 5627
rect 1869 5593 1903 5627
rect 1903 5593 1912 5627
rect 1860 5584 1912 5593
rect 46572 5516 46624 5568
rect 30398 5414 30450 5466
rect 30462 5414 30514 5466
rect 30526 5414 30578 5466
rect 30590 5414 30642 5466
rect 30654 5414 30706 5466
rect 59846 5414 59898 5466
rect 59910 5414 59962 5466
rect 59974 5414 60026 5466
rect 60038 5414 60090 5466
rect 60102 5414 60154 5466
rect 89294 5414 89346 5466
rect 89358 5414 89410 5466
rect 89422 5414 89474 5466
rect 89486 5414 89538 5466
rect 89550 5414 89602 5466
rect 83004 5287 83056 5296
rect 83004 5253 83013 5287
rect 83013 5253 83047 5287
rect 83047 5253 83056 5287
rect 83004 5244 83056 5253
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 82820 5219 82872 5228
rect 82820 5185 82829 5219
rect 82829 5185 82863 5219
rect 82863 5185 82872 5219
rect 82820 5176 82872 5185
rect 115664 5176 115716 5228
rect 61016 4972 61068 5024
rect 117964 5015 118016 5024
rect 117964 4981 117973 5015
rect 117973 4981 118007 5015
rect 118007 4981 118016 5015
rect 117964 4972 118016 4981
rect 15674 4870 15726 4922
rect 15738 4870 15790 4922
rect 15802 4870 15854 4922
rect 15866 4870 15918 4922
rect 15930 4870 15982 4922
rect 45122 4870 45174 4922
rect 45186 4870 45238 4922
rect 45250 4870 45302 4922
rect 45314 4870 45366 4922
rect 45378 4870 45430 4922
rect 74570 4870 74622 4922
rect 74634 4870 74686 4922
rect 74698 4870 74750 4922
rect 74762 4870 74814 4922
rect 74826 4870 74878 4922
rect 104018 4870 104070 4922
rect 104082 4870 104134 4922
rect 104146 4870 104198 4922
rect 104210 4870 104262 4922
rect 104274 4870 104326 4922
rect 42616 4564 42668 4616
rect 79232 4564 79284 4616
rect 37648 4428 37700 4480
rect 70584 4428 70636 4480
rect 71412 4428 71464 4480
rect 115664 4496 115716 4548
rect 117780 4539 117832 4548
rect 117780 4505 117789 4539
rect 117789 4505 117823 4539
rect 117823 4505 117832 4539
rect 117780 4496 117832 4505
rect 30398 4326 30450 4378
rect 30462 4326 30514 4378
rect 30526 4326 30578 4378
rect 30590 4326 30642 4378
rect 30654 4326 30706 4378
rect 59846 4326 59898 4378
rect 59910 4326 59962 4378
rect 59974 4326 60026 4378
rect 60038 4326 60090 4378
rect 60102 4326 60154 4378
rect 89294 4326 89346 4378
rect 89358 4326 89410 4378
rect 89422 4326 89474 4378
rect 89486 4326 89538 4378
rect 89550 4326 89602 4378
rect 82636 4267 82688 4276
rect 1400 4088 1452 4140
rect 1768 4088 1820 4140
rect 2596 4088 2648 4140
rect 35716 4088 35768 4140
rect 59268 4088 59320 4140
rect 59636 4088 59688 4140
rect 59820 4088 59872 4140
rect 61752 4156 61804 4208
rect 82636 4233 82645 4267
rect 82645 4233 82679 4267
rect 82679 4233 82688 4267
rect 82636 4224 82688 4233
rect 73068 4156 73120 4208
rect 85488 4156 85540 4208
rect 119804 4156 119856 4208
rect 1952 4020 2004 4072
rect 57244 4020 57296 4072
rect 57336 4020 57388 4072
rect 65064 4020 65116 4072
rect 72608 4020 72660 4072
rect 77208 4088 77260 4140
rect 79232 4131 79284 4140
rect 79232 4097 79241 4131
rect 79241 4097 79275 4131
rect 79275 4097 79284 4131
rect 79232 4088 79284 4097
rect 107476 4088 107528 4140
rect 116860 4131 116912 4140
rect 116860 4097 116869 4131
rect 116869 4097 116903 4131
rect 116903 4097 116912 4131
rect 116860 4088 116912 4097
rect 1492 3952 1544 4004
rect 2136 3952 2188 4004
rect 31484 3884 31536 3936
rect 57336 3884 57388 3936
rect 74172 3952 74224 4004
rect 59360 3927 59412 3936
rect 59360 3893 59369 3927
rect 59369 3893 59403 3927
rect 59403 3893 59412 3927
rect 59360 3884 59412 3893
rect 59636 3884 59688 3936
rect 61752 3884 61804 3936
rect 73068 3884 73120 3936
rect 73160 3884 73212 3936
rect 73712 3884 73764 3936
rect 74080 3884 74132 3936
rect 82728 4063 82780 4072
rect 82728 4029 82737 4063
rect 82737 4029 82771 4063
rect 82771 4029 82780 4063
rect 82728 4020 82780 4029
rect 74356 3952 74408 4004
rect 82636 3952 82688 4004
rect 77024 3884 77076 3936
rect 79508 3884 79560 3936
rect 82820 3884 82872 3936
rect 117964 3884 118016 3936
rect 118056 3927 118108 3936
rect 118056 3893 118065 3927
rect 118065 3893 118099 3927
rect 118099 3893 118108 3927
rect 118056 3884 118108 3893
rect 15674 3782 15726 3834
rect 15738 3782 15790 3834
rect 15802 3782 15854 3834
rect 15866 3782 15918 3834
rect 15930 3782 15982 3834
rect 45122 3782 45174 3834
rect 45186 3782 45238 3834
rect 45250 3782 45302 3834
rect 45314 3782 45366 3834
rect 45378 3782 45430 3834
rect 74570 3782 74622 3834
rect 74634 3782 74686 3834
rect 74698 3782 74750 3834
rect 74762 3782 74814 3834
rect 74826 3782 74878 3834
rect 104018 3782 104070 3834
rect 104082 3782 104134 3834
rect 104146 3782 104198 3834
rect 104210 3782 104262 3834
rect 104274 3782 104326 3834
rect 5448 3680 5500 3732
rect 45652 3680 45704 3732
rect 20720 3544 20772 3596
rect 40132 3612 40184 3664
rect 56968 3680 57020 3732
rect 57060 3680 57112 3732
rect 59636 3723 59688 3732
rect 33600 3544 33652 3596
rect 57980 3612 58032 3664
rect 59636 3689 59645 3723
rect 59645 3689 59679 3723
rect 59679 3689 59688 3723
rect 59636 3680 59688 3689
rect 72332 3680 72384 3732
rect 117136 3680 117188 3732
rect 59820 3612 59872 3664
rect 61016 3612 61068 3664
rect 72240 3612 72292 3664
rect 73068 3612 73120 3664
rect 74080 3612 74132 3664
rect 117688 3680 117740 3732
rect 46848 3544 46900 3596
rect 57060 3544 57112 3596
rect 57152 3544 57204 3596
rect 58072 3544 58124 3596
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 664 3408 716 3460
rect 32128 3476 32180 3528
rect 33784 3476 33836 3528
rect 40316 3476 40368 3528
rect 40592 3476 40644 3528
rect 41512 3476 41564 3528
rect 42432 3476 42484 3528
rect 34980 3408 35032 3460
rect 40408 3408 40460 3460
rect 45744 3476 45796 3528
rect 47216 3476 47268 3528
rect 47952 3476 48004 3528
rect 48044 3476 48096 3528
rect 50712 3476 50764 3528
rect 47308 3408 47360 3460
rect 52184 3476 52236 3528
rect 57612 3519 57664 3528
rect 57612 3485 57621 3519
rect 57621 3485 57655 3519
rect 57655 3485 57664 3519
rect 57612 3476 57664 3485
rect 61660 3544 61712 3596
rect 97816 3544 97868 3596
rect 58256 3515 58308 3528
rect 58256 3481 58257 3515
rect 58257 3481 58291 3515
rect 58291 3481 58308 3515
rect 58256 3476 58308 3481
rect 58532 3476 58584 3528
rect 68468 3476 68520 3528
rect 70768 3476 70820 3528
rect 71596 3519 71648 3528
rect 71596 3485 71605 3519
rect 71605 3485 71639 3519
rect 71639 3485 71648 3519
rect 71596 3476 71648 3485
rect 72148 3476 72200 3528
rect 73160 3476 73212 3528
rect 74172 3519 74224 3528
rect 74172 3485 74181 3519
rect 74181 3485 74215 3519
rect 74215 3485 74224 3519
rect 74172 3476 74224 3485
rect 74908 3476 74960 3528
rect 78036 3476 78088 3528
rect 59544 3451 59596 3460
rect 59544 3417 59553 3451
rect 59553 3417 59587 3451
rect 59587 3417 59596 3451
rect 59544 3408 59596 3417
rect 60280 3408 60332 3460
rect 66996 3408 67048 3460
rect 101496 3408 101548 3460
rect 1308 3340 1360 3392
rect 2872 3340 2924 3392
rect 41788 3340 41840 3392
rect 42432 3340 42484 3392
rect 42800 3340 42852 3392
rect 45836 3383 45888 3392
rect 45836 3349 45845 3383
rect 45845 3349 45879 3383
rect 45879 3349 45888 3383
rect 45836 3340 45888 3349
rect 46848 3383 46900 3392
rect 46848 3349 46857 3383
rect 46857 3349 46891 3383
rect 46891 3349 46900 3383
rect 46848 3340 46900 3349
rect 47492 3383 47544 3392
rect 47492 3349 47501 3383
rect 47501 3349 47535 3383
rect 47535 3349 47544 3383
rect 47492 3340 47544 3349
rect 47584 3340 47636 3392
rect 50804 3340 50856 3392
rect 50896 3340 50948 3392
rect 57152 3340 57204 3392
rect 57336 3340 57388 3392
rect 58164 3340 58216 3392
rect 70216 3340 70268 3392
rect 70860 3340 70912 3392
rect 72056 3383 72108 3392
rect 72056 3349 72065 3383
rect 72065 3349 72099 3383
rect 72099 3349 72108 3383
rect 72056 3340 72108 3349
rect 74172 3340 74224 3392
rect 74540 3340 74592 3392
rect 75460 3340 75512 3392
rect 76012 3340 76064 3392
rect 77116 3340 77168 3392
rect 77484 3340 77536 3392
rect 117412 3519 117464 3528
rect 116676 3340 116728 3392
rect 117412 3485 117421 3519
rect 117421 3485 117455 3519
rect 117455 3485 117464 3519
rect 117412 3476 117464 3485
rect 117872 3519 117924 3528
rect 117872 3485 117881 3519
rect 117881 3485 117915 3519
rect 117915 3485 117924 3519
rect 117872 3476 117924 3485
rect 30398 3238 30450 3290
rect 30462 3238 30514 3290
rect 30526 3238 30578 3290
rect 30590 3238 30642 3290
rect 30654 3238 30706 3290
rect 59846 3238 59898 3290
rect 59910 3238 59962 3290
rect 59974 3238 60026 3290
rect 60038 3238 60090 3290
rect 60102 3238 60154 3290
rect 89294 3238 89346 3290
rect 89358 3238 89410 3290
rect 89422 3238 89474 3290
rect 89486 3238 89538 3290
rect 89550 3238 89602 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 2596 3136 2648 3188
rect 2780 3068 2832 3120
rect 10232 3136 10284 3188
rect 20720 3179 20772 3188
rect 20720 3145 20729 3179
rect 20729 3145 20763 3179
rect 20763 3145 20772 3179
rect 20720 3136 20772 3145
rect 24492 3136 24544 3188
rect 28908 3179 28960 3188
rect 2596 3000 2648 3052
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 7196 3000 7248 3052
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 12348 3000 12400 3052
rect 14188 3000 14240 3052
rect 20628 3000 20680 3052
rect 23112 3000 23164 3052
rect 24492 3043 24544 3052
rect 24492 3009 24501 3043
rect 24501 3009 24535 3043
rect 24535 3009 24544 3043
rect 24492 3000 24544 3009
rect 27620 3043 27672 3052
rect 27620 3009 27629 3043
rect 27629 3009 27663 3043
rect 27663 3009 27672 3043
rect 27620 3000 27672 3009
rect 7748 2932 7800 2984
rect 28908 3145 28917 3179
rect 28917 3145 28951 3179
rect 28951 3145 28960 3179
rect 28908 3136 28960 3145
rect 29644 3179 29696 3188
rect 29644 3145 29653 3179
rect 29653 3145 29687 3179
rect 29687 3145 29696 3179
rect 29644 3136 29696 3145
rect 41236 3136 41288 3188
rect 32956 3111 33008 3120
rect 32956 3077 32965 3111
rect 32965 3077 32999 3111
rect 32999 3077 33008 3111
rect 32956 3068 33008 3077
rect 28908 3000 28960 3052
rect 20 2864 72 2916
rect 5172 2796 5224 2848
rect 5816 2796 5868 2848
rect 7104 2796 7156 2848
rect 12624 2796 12676 2848
rect 24768 2796 24820 2848
rect 26424 2839 26476 2848
rect 26424 2805 26433 2839
rect 26433 2805 26467 2839
rect 26467 2805 26476 2839
rect 26424 2796 26476 2805
rect 33600 3043 33652 3052
rect 33600 3009 33609 3043
rect 33609 3009 33643 3043
rect 33643 3009 33652 3043
rect 33600 3000 33652 3009
rect 34796 3000 34848 3052
rect 35440 3000 35492 3052
rect 36084 3000 36136 3052
rect 37648 3043 37700 3052
rect 37648 3009 37657 3043
rect 37657 3009 37691 3043
rect 37691 3009 37700 3043
rect 37648 3000 37700 3009
rect 37740 2975 37792 2984
rect 37740 2941 37749 2975
rect 37749 2941 37783 2975
rect 37783 2941 37792 2975
rect 37740 2932 37792 2941
rect 37832 2975 37884 2984
rect 37832 2941 37841 2975
rect 37841 2941 37875 2975
rect 37875 2941 37884 2975
rect 37832 2932 37884 2941
rect 35716 2907 35768 2916
rect 35716 2873 35725 2907
rect 35725 2873 35759 2907
rect 35759 2873 35768 2907
rect 35716 2864 35768 2873
rect 41788 3136 41840 3188
rect 42800 3136 42852 3188
rect 42984 3111 43036 3120
rect 42984 3077 42993 3111
rect 42993 3077 43027 3111
rect 43027 3077 43036 3111
rect 47676 3136 47728 3188
rect 42984 3068 43036 3077
rect 39580 3043 39632 3052
rect 39580 3009 39589 3043
rect 39589 3009 39623 3043
rect 39623 3009 39632 3043
rect 39580 3000 39632 3009
rect 40408 3043 40460 3052
rect 40408 3009 40417 3043
rect 40417 3009 40451 3043
rect 40451 3009 40460 3043
rect 40408 3000 40460 3009
rect 41696 3000 41748 3052
rect 41972 3000 42024 3052
rect 43812 3000 43864 3052
rect 45376 3043 45428 3052
rect 45376 3009 45385 3043
rect 45385 3009 45419 3043
rect 45419 3009 45428 3043
rect 45376 3000 45428 3009
rect 46388 3000 46440 3052
rect 47124 3068 47176 3120
rect 47860 3136 47912 3188
rect 57612 3136 57664 3188
rect 58072 3179 58124 3188
rect 58072 3145 58081 3179
rect 58081 3145 58115 3179
rect 58115 3145 58124 3179
rect 58072 3136 58124 3145
rect 47584 3000 47636 3052
rect 47952 3043 48004 3052
rect 47952 3009 47961 3043
rect 47961 3009 47995 3043
rect 47995 3009 48004 3043
rect 47952 3000 48004 3009
rect 40224 2932 40276 2984
rect 40684 2975 40736 2984
rect 40684 2941 40693 2975
rect 40693 2941 40727 2975
rect 40727 2941 40736 2975
rect 40684 2932 40736 2941
rect 43260 2975 43312 2984
rect 43260 2941 43269 2975
rect 43269 2941 43303 2975
rect 43303 2941 43312 2975
rect 43260 2932 43312 2941
rect 45836 2932 45888 2984
rect 51172 3043 51224 3052
rect 51172 3009 51181 3043
rect 51181 3009 51215 3043
rect 51215 3009 51224 3043
rect 51172 3000 51224 3009
rect 52736 3000 52788 3052
rect 52828 3000 52880 3052
rect 54116 3068 54168 3120
rect 56692 3068 56744 3120
rect 56968 3111 57020 3120
rect 56968 3077 56977 3111
rect 56977 3077 57011 3111
rect 57011 3077 57020 3111
rect 56968 3068 57020 3077
rect 57152 3068 57204 3120
rect 57980 3068 58032 3120
rect 76012 3136 76064 3188
rect 59544 3068 59596 3120
rect 61660 3068 61712 3120
rect 61752 3068 61804 3120
rect 70308 3068 70360 3120
rect 70584 3111 70636 3120
rect 70584 3077 70593 3111
rect 70593 3077 70627 3111
rect 70627 3077 70636 3111
rect 70584 3068 70636 3077
rect 74540 3111 74592 3120
rect 74540 3077 74549 3111
rect 74549 3077 74583 3111
rect 74583 3077 74592 3111
rect 74540 3068 74592 3077
rect 75368 3068 75420 3120
rect 77116 3136 77168 3188
rect 85304 3136 85356 3188
rect 77024 3068 77076 3120
rect 102784 3136 102836 3188
rect 104256 3136 104308 3188
rect 117136 3179 117188 3188
rect 103980 3068 104032 3120
rect 107476 3111 107528 3120
rect 107476 3077 107485 3111
rect 107485 3077 107519 3111
rect 107519 3077 107528 3111
rect 107476 3068 107528 3077
rect 109776 3068 109828 3120
rect 55588 3000 55640 3052
rect 57704 3000 57756 3052
rect 50620 2932 50672 2984
rect 48044 2864 48096 2916
rect 28356 2796 28408 2848
rect 31576 2796 31628 2848
rect 32864 2796 32916 2848
rect 36268 2839 36320 2848
rect 36268 2805 36277 2839
rect 36277 2805 36311 2839
rect 36311 2805 36320 2839
rect 36268 2796 36320 2805
rect 37648 2796 37700 2848
rect 39396 2839 39448 2848
rect 39396 2805 39405 2839
rect 39405 2805 39439 2839
rect 39439 2805 39448 2839
rect 39396 2796 39448 2805
rect 40040 2839 40092 2848
rect 40040 2805 40049 2839
rect 40049 2805 40083 2839
rect 40083 2805 40092 2839
rect 40040 2796 40092 2805
rect 42616 2839 42668 2848
rect 42616 2805 42625 2839
rect 42625 2805 42659 2839
rect 42659 2805 42668 2839
rect 42616 2796 42668 2805
rect 46204 2839 46256 2848
rect 46204 2805 46213 2839
rect 46213 2805 46247 2839
rect 46247 2805 46256 2839
rect 46204 2796 46256 2805
rect 46296 2796 46348 2848
rect 57428 2932 57480 2984
rect 59728 3043 59780 3052
rect 57980 2932 58032 2984
rect 59452 2975 59504 2984
rect 59452 2941 59461 2975
rect 59461 2941 59495 2975
rect 59495 2941 59504 2975
rect 59452 2932 59504 2941
rect 59728 3009 59737 3043
rect 59737 3009 59771 3043
rect 59771 3009 59780 3043
rect 59728 3000 59780 3009
rect 61844 3000 61896 3052
rect 64052 3000 64104 3052
rect 64512 3000 64564 3052
rect 66720 3000 66772 3052
rect 66996 3043 67048 3052
rect 66996 3009 67005 3043
rect 67005 3009 67039 3043
rect 67039 3009 67048 3043
rect 66996 3000 67048 3009
rect 68284 3000 68336 3052
rect 69572 3000 69624 3052
rect 70400 3043 70452 3052
rect 70400 3009 70409 3043
rect 70409 3009 70443 3043
rect 70443 3009 70452 3043
rect 70400 3000 70452 3009
rect 60004 2932 60056 2984
rect 69940 2932 69992 2984
rect 71320 3000 71372 3052
rect 72240 3043 72292 3052
rect 72240 3009 72249 3043
rect 72249 3009 72283 3043
rect 72283 3009 72292 3043
rect 72240 3000 72292 3009
rect 72332 3043 72384 3052
rect 72332 3009 72341 3043
rect 72341 3009 72375 3043
rect 72375 3009 72384 3043
rect 72332 3000 72384 3009
rect 64604 2907 64656 2916
rect 48320 2796 48372 2848
rect 50896 2796 50948 2848
rect 52920 2839 52972 2848
rect 52920 2805 52929 2839
rect 52929 2805 52963 2839
rect 52963 2805 52972 2839
rect 52920 2796 52972 2805
rect 55404 2796 55456 2848
rect 55864 2796 55916 2848
rect 56692 2796 56744 2848
rect 57980 2796 58032 2848
rect 58072 2796 58124 2848
rect 58256 2796 58308 2848
rect 58808 2839 58860 2848
rect 58808 2805 58817 2839
rect 58817 2805 58851 2839
rect 58851 2805 58860 2839
rect 58808 2796 58860 2805
rect 64604 2873 64613 2907
rect 64613 2873 64647 2907
rect 64647 2873 64656 2907
rect 64604 2864 64656 2873
rect 66168 2907 66220 2916
rect 66168 2873 66177 2907
rect 66177 2873 66211 2907
rect 66211 2873 66220 2907
rect 66168 2864 66220 2873
rect 68468 2864 68520 2916
rect 61752 2796 61804 2848
rect 61936 2839 61988 2848
rect 61936 2805 61945 2839
rect 61945 2805 61979 2839
rect 61979 2805 61988 2839
rect 61936 2796 61988 2805
rect 63500 2796 63552 2848
rect 66352 2796 66404 2848
rect 68100 2796 68152 2848
rect 69664 2839 69716 2848
rect 69664 2805 69673 2839
rect 69673 2805 69707 2839
rect 69707 2805 69716 2839
rect 69664 2796 69716 2805
rect 71228 2864 71280 2916
rect 72332 2864 72384 2916
rect 76840 3043 76892 3052
rect 76840 3009 76849 3043
rect 76849 3009 76883 3043
rect 76883 3009 76892 3043
rect 76840 3000 76892 3009
rect 77300 3000 77352 3052
rect 80704 3000 80756 3052
rect 87236 3043 87288 3052
rect 87236 3009 87245 3043
rect 87245 3009 87279 3043
rect 87279 3009 87288 3043
rect 87236 3000 87288 3009
rect 101496 3043 101548 3052
rect 101496 3009 101505 3043
rect 101505 3009 101539 3043
rect 101539 3009 101548 3043
rect 101496 3000 101548 3009
rect 102692 3043 102744 3052
rect 102692 3009 102701 3043
rect 102701 3009 102735 3043
rect 102735 3009 102744 3043
rect 102692 3000 102744 3009
rect 102784 3000 102836 3052
rect 110236 3000 110288 3052
rect 111432 3000 111484 3052
rect 116216 3043 116268 3052
rect 116216 3009 116225 3043
rect 116225 3009 116259 3043
rect 116259 3009 116268 3043
rect 116216 3000 116268 3009
rect 117136 3145 117145 3179
rect 117145 3145 117179 3179
rect 117179 3145 117188 3179
rect 117136 3136 117188 3145
rect 118516 3068 118568 3120
rect 117412 3000 117464 3052
rect 117780 3043 117832 3052
rect 117780 3009 117789 3043
rect 117789 3009 117823 3043
rect 117823 3009 117832 3043
rect 117780 3000 117832 3009
rect 75092 2864 75144 2916
rect 75736 2864 75788 2916
rect 76472 2907 76524 2916
rect 76472 2873 76481 2907
rect 76481 2873 76515 2907
rect 76515 2873 76524 2907
rect 76472 2864 76524 2873
rect 73436 2796 73488 2848
rect 75552 2796 75604 2848
rect 76932 2932 76984 2984
rect 77116 2932 77168 2984
rect 76840 2864 76892 2916
rect 89168 2864 89220 2916
rect 107660 2907 107712 2916
rect 107660 2873 107669 2907
rect 107669 2873 107703 2907
rect 107703 2873 107712 2907
rect 107660 2864 107712 2873
rect 109500 2864 109552 2916
rect 110236 2864 110288 2916
rect 81164 2796 81216 2848
rect 86960 2796 87012 2848
rect 98552 2796 98604 2848
rect 102416 2796 102468 2848
rect 109776 2839 109828 2848
rect 109776 2805 109785 2839
rect 109785 2805 109819 2839
rect 109819 2805 109828 2839
rect 109776 2796 109828 2805
rect 115940 2796 115992 2848
rect 15674 2694 15726 2746
rect 15738 2694 15790 2746
rect 15802 2694 15854 2746
rect 15866 2694 15918 2746
rect 15930 2694 15982 2746
rect 45122 2694 45174 2746
rect 45186 2694 45238 2746
rect 45250 2694 45302 2746
rect 45314 2694 45366 2746
rect 45378 2694 45430 2746
rect 74570 2694 74622 2746
rect 74634 2694 74686 2746
rect 74698 2694 74750 2746
rect 74762 2694 74814 2746
rect 74826 2694 74878 2746
rect 104018 2694 104070 2746
rect 104082 2694 104134 2746
rect 104146 2694 104198 2746
rect 104210 2694 104262 2746
rect 104274 2694 104326 2746
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 14648 2635 14700 2644
rect 14648 2601 14657 2635
rect 14657 2601 14691 2635
rect 14691 2601 14700 2635
rect 14648 2592 14700 2601
rect 19432 2592 19484 2644
rect 22468 2592 22520 2644
rect 23112 2592 23164 2644
rect 23296 2635 23348 2644
rect 23296 2601 23305 2635
rect 23305 2601 23339 2635
rect 23339 2601 23348 2635
rect 23296 2592 23348 2601
rect 25412 2635 25464 2644
rect 25412 2601 25421 2635
rect 25421 2601 25455 2635
rect 25455 2601 25464 2635
rect 25412 2592 25464 2601
rect 27620 2592 27672 2644
rect 28816 2635 28868 2644
rect 28816 2601 28825 2635
rect 28825 2601 28859 2635
rect 28859 2601 28868 2635
rect 28816 2592 28868 2601
rect 32128 2635 32180 2644
rect 32128 2601 32137 2635
rect 32137 2601 32171 2635
rect 32171 2601 32180 2635
rect 32128 2592 32180 2601
rect 9680 2524 9732 2576
rect 58716 2592 58768 2644
rect 59452 2592 59504 2644
rect 38016 2524 38068 2576
rect 38568 2524 38620 2576
rect 40224 2524 40276 2576
rect 40684 2524 40736 2576
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 3240 2388 3292 2440
rect 4528 2388 4580 2440
rect 9036 2388 9088 2440
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 11612 2388 11664 2440
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 10968 2320 11020 2372
rect 13544 2320 13596 2372
rect 16120 2456 16172 2508
rect 27528 2499 27580 2508
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 17408 2388 17460 2440
rect 19432 2431 19484 2440
rect 18236 2320 18288 2372
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19984 2388 20036 2440
rect 19708 2320 19760 2372
rect 21916 2388 21968 2440
rect 22560 2388 22612 2440
rect 23204 2388 23256 2440
rect 24676 2388 24728 2440
rect 24860 2388 24912 2440
rect 25136 2388 25188 2440
rect 27068 2388 27120 2440
rect 27528 2465 27537 2499
rect 27537 2465 27571 2499
rect 27571 2465 27580 2499
rect 27528 2456 27580 2465
rect 27712 2388 27764 2440
rect 29736 2456 29788 2508
rect 29828 2456 29880 2508
rect 32772 2499 32824 2508
rect 28816 2388 28868 2440
rect 29000 2431 29052 2440
rect 29000 2397 29009 2431
rect 29009 2397 29043 2431
rect 29043 2397 29052 2431
rect 29000 2388 29052 2397
rect 29644 2388 29696 2440
rect 30932 2431 30984 2440
rect 30932 2397 30941 2431
rect 30941 2397 30975 2431
rect 30975 2397 30984 2431
rect 30932 2388 30984 2397
rect 31576 2431 31628 2440
rect 31576 2397 31585 2431
rect 31585 2397 31619 2431
rect 31619 2397 31628 2431
rect 31576 2388 31628 2397
rect 28264 2320 28316 2372
rect 32772 2465 32781 2499
rect 32781 2465 32815 2499
rect 32815 2465 32824 2499
rect 32772 2456 32824 2465
rect 34704 2499 34756 2508
rect 7012 2295 7064 2304
rect 7012 2261 7021 2295
rect 7021 2261 7055 2295
rect 7055 2261 7064 2295
rect 7012 2252 7064 2261
rect 10140 2295 10192 2304
rect 10140 2261 10149 2295
rect 10149 2261 10183 2295
rect 10183 2261 10192 2295
rect 10140 2252 10192 2261
rect 12256 2252 12308 2304
rect 15476 2252 15528 2304
rect 16120 2252 16172 2304
rect 17500 2295 17552 2304
rect 17500 2261 17509 2295
rect 17509 2261 17543 2295
rect 17543 2261 17552 2295
rect 17500 2252 17552 2261
rect 18052 2252 18104 2304
rect 18696 2252 18748 2304
rect 24492 2252 24544 2304
rect 24676 2252 24728 2304
rect 26148 2252 26200 2304
rect 27160 2252 27212 2304
rect 27344 2252 27396 2304
rect 28172 2295 28224 2304
rect 28172 2261 28181 2295
rect 28181 2261 28215 2295
rect 28215 2261 28224 2295
rect 28172 2252 28224 2261
rect 29736 2295 29788 2304
rect 29736 2261 29745 2295
rect 29745 2261 29779 2295
rect 29779 2261 29788 2295
rect 29736 2252 29788 2261
rect 30748 2295 30800 2304
rect 30748 2261 30757 2295
rect 30757 2261 30791 2295
rect 30791 2261 30800 2295
rect 30748 2252 30800 2261
rect 31300 2252 31352 2304
rect 31668 2252 31720 2304
rect 34704 2465 34713 2499
rect 34713 2465 34747 2499
rect 34747 2465 34756 2499
rect 34704 2456 34756 2465
rect 37832 2456 37884 2508
rect 45560 2524 45612 2576
rect 47584 2567 47636 2576
rect 47584 2533 47593 2567
rect 47593 2533 47627 2567
rect 47627 2533 47636 2567
rect 47584 2524 47636 2533
rect 42616 2456 42668 2508
rect 46756 2499 46808 2508
rect 46756 2465 46765 2499
rect 46765 2465 46799 2499
rect 46799 2465 46808 2499
rect 46756 2456 46808 2465
rect 48044 2499 48096 2508
rect 48044 2465 48053 2499
rect 48053 2465 48087 2499
rect 48087 2465 48096 2499
rect 48044 2456 48096 2465
rect 50436 2524 50488 2576
rect 50804 2524 50856 2576
rect 52736 2567 52788 2576
rect 52000 2499 52052 2508
rect 33508 2252 33560 2304
rect 34704 2252 34756 2304
rect 36268 2388 36320 2440
rect 37648 2431 37700 2440
rect 37648 2397 37657 2431
rect 37657 2397 37691 2431
rect 37691 2397 37700 2431
rect 37648 2388 37700 2397
rect 38660 2431 38712 2440
rect 38660 2397 38669 2431
rect 38669 2397 38703 2431
rect 38703 2397 38712 2431
rect 38660 2388 38712 2397
rect 39304 2431 39356 2440
rect 39304 2397 39313 2431
rect 39313 2397 39347 2431
rect 39347 2397 39356 2431
rect 39304 2388 39356 2397
rect 40132 2388 40184 2440
rect 42708 2431 42760 2440
rect 42708 2397 42717 2431
rect 42717 2397 42751 2431
rect 42751 2397 42760 2431
rect 42708 2388 42760 2397
rect 45928 2388 45980 2440
rect 36544 2320 36596 2372
rect 39856 2320 39908 2372
rect 37372 2252 37424 2304
rect 39948 2252 40000 2304
rect 41788 2363 41840 2372
rect 41788 2329 41797 2363
rect 41797 2329 41831 2363
rect 41831 2329 41840 2363
rect 41788 2320 41840 2329
rect 40500 2252 40552 2304
rect 44456 2252 44508 2304
rect 45560 2295 45612 2304
rect 45560 2261 45569 2295
rect 45569 2261 45603 2295
rect 45603 2261 45612 2295
rect 49148 2388 49200 2440
rect 52000 2465 52009 2499
rect 52009 2465 52043 2499
rect 52043 2465 52052 2499
rect 52000 2456 52052 2465
rect 52736 2533 52745 2567
rect 52745 2533 52779 2567
rect 52779 2533 52788 2567
rect 52736 2524 52788 2533
rect 52920 2456 52972 2508
rect 54024 2524 54076 2576
rect 62764 2592 62816 2644
rect 63776 2592 63828 2644
rect 66720 2635 66772 2644
rect 66720 2601 66729 2635
rect 66729 2601 66763 2635
rect 66763 2601 66772 2635
rect 66720 2592 66772 2601
rect 70768 2635 70820 2644
rect 60004 2524 60056 2576
rect 56416 2456 56468 2508
rect 56784 2499 56836 2508
rect 56784 2465 56793 2499
rect 56793 2465 56827 2499
rect 56827 2465 56836 2499
rect 56784 2456 56836 2465
rect 57796 2456 57848 2508
rect 62580 2524 62632 2576
rect 46756 2320 46808 2372
rect 45560 2252 45612 2261
rect 46664 2295 46716 2304
rect 46664 2261 46673 2295
rect 46673 2261 46707 2295
rect 46707 2261 46716 2295
rect 46664 2252 46716 2261
rect 47952 2295 48004 2304
rect 47952 2261 47961 2295
rect 47961 2261 47995 2295
rect 47995 2261 48004 2295
rect 47952 2252 48004 2261
rect 48964 2252 49016 2304
rect 50252 2252 50304 2304
rect 53932 2388 53984 2440
rect 54116 2431 54168 2440
rect 54116 2397 54125 2431
rect 54125 2397 54159 2431
rect 54159 2397 54168 2431
rect 54116 2388 54168 2397
rect 54760 2431 54812 2440
rect 54760 2397 54769 2431
rect 54769 2397 54803 2431
rect 54803 2397 54812 2431
rect 54760 2388 54812 2397
rect 51632 2320 51684 2372
rect 54024 2320 54076 2372
rect 55864 2363 55916 2372
rect 55864 2329 55873 2363
rect 55873 2329 55907 2363
rect 55907 2329 55916 2363
rect 55864 2320 55916 2329
rect 56692 2388 56744 2440
rect 58164 2431 58216 2440
rect 58164 2397 58173 2431
rect 58173 2397 58207 2431
rect 58207 2397 58216 2431
rect 58164 2388 58216 2397
rect 61292 2388 61344 2440
rect 61476 2388 61528 2440
rect 63408 2431 63460 2440
rect 63408 2397 63417 2431
rect 63417 2397 63451 2431
rect 63451 2397 63460 2431
rect 63408 2388 63460 2397
rect 64052 2431 64104 2440
rect 64052 2397 64061 2431
rect 64061 2397 64095 2431
rect 64095 2397 64104 2431
rect 64052 2388 64104 2397
rect 65984 2431 66036 2440
rect 59360 2320 59412 2372
rect 65984 2397 65993 2431
rect 65993 2397 66027 2431
rect 66027 2397 66036 2431
rect 65984 2388 66036 2397
rect 66076 2388 66128 2440
rect 67456 2524 67508 2576
rect 68928 2567 68980 2576
rect 68928 2533 68937 2567
rect 68937 2533 68971 2567
rect 68971 2533 68980 2567
rect 68928 2524 68980 2533
rect 70400 2524 70452 2576
rect 70768 2601 70777 2635
rect 70777 2601 70811 2635
rect 70811 2601 70820 2635
rect 70768 2592 70820 2601
rect 71320 2592 71372 2644
rect 72332 2592 72384 2644
rect 82452 2592 82504 2644
rect 82544 2635 82596 2644
rect 82544 2601 82553 2635
rect 82553 2601 82587 2635
rect 82587 2601 82596 2635
rect 82544 2592 82596 2601
rect 82728 2592 82780 2644
rect 102232 2635 102284 2644
rect 102232 2601 102241 2635
rect 102241 2601 102275 2635
rect 102275 2601 102284 2635
rect 102232 2592 102284 2601
rect 103336 2635 103388 2644
rect 103336 2601 103345 2635
rect 103345 2601 103379 2635
rect 103379 2601 103388 2635
rect 103336 2592 103388 2601
rect 104532 2592 104584 2644
rect 114744 2592 114796 2644
rect 67364 2388 67416 2440
rect 69664 2431 69716 2440
rect 69664 2397 69673 2431
rect 69673 2397 69707 2431
rect 69707 2397 69716 2431
rect 69664 2388 69716 2397
rect 69940 2456 69992 2508
rect 71872 2456 71924 2508
rect 72056 2499 72108 2508
rect 72056 2465 72065 2499
rect 72065 2465 72099 2499
rect 72099 2465 72108 2499
rect 72056 2456 72108 2465
rect 70584 2388 70636 2440
rect 71228 2388 71280 2440
rect 71320 2388 71372 2440
rect 73528 2456 73580 2508
rect 73988 2499 74040 2508
rect 73988 2465 73997 2499
rect 73997 2465 74031 2499
rect 74031 2465 74040 2499
rect 73988 2456 74040 2465
rect 77024 2456 77076 2508
rect 77208 2456 77260 2508
rect 118240 2524 118292 2576
rect 73712 2388 73764 2440
rect 51816 2295 51868 2304
rect 51816 2261 51825 2295
rect 51825 2261 51859 2295
rect 51859 2261 51868 2295
rect 51816 2252 51868 2261
rect 51908 2295 51960 2304
rect 51908 2261 51917 2295
rect 51917 2261 51951 2295
rect 51951 2261 51960 2295
rect 53104 2295 53156 2304
rect 51908 2252 51960 2261
rect 53104 2261 53113 2295
rect 53113 2261 53147 2295
rect 53147 2261 53156 2295
rect 53104 2252 53156 2261
rect 53472 2252 53524 2304
rect 55956 2295 56008 2304
rect 55956 2261 55965 2295
rect 55965 2261 55999 2295
rect 55999 2261 56008 2295
rect 55956 2252 56008 2261
rect 58256 2295 58308 2304
rect 58256 2261 58265 2295
rect 58265 2261 58299 2295
rect 58299 2261 58308 2295
rect 58256 2252 58308 2261
rect 61016 2295 61068 2304
rect 61016 2261 61025 2295
rect 61025 2261 61059 2295
rect 61059 2261 61068 2295
rect 61016 2252 61068 2261
rect 63132 2252 63184 2304
rect 66812 2320 66864 2372
rect 67272 2320 67324 2372
rect 71044 2320 71096 2372
rect 71136 2320 71188 2372
rect 65708 2252 65760 2304
rect 67180 2295 67232 2304
rect 67180 2261 67189 2295
rect 67189 2261 67223 2295
rect 67223 2261 67232 2295
rect 67180 2252 67232 2261
rect 67640 2252 67692 2304
rect 68928 2252 68980 2304
rect 73620 2295 73672 2304
rect 73620 2261 73629 2295
rect 73629 2261 73663 2295
rect 73663 2261 73672 2295
rect 73620 2252 73672 2261
rect 74632 2295 74684 2304
rect 74632 2261 74641 2295
rect 74641 2261 74675 2295
rect 74675 2261 74684 2295
rect 74632 2252 74684 2261
rect 75828 2388 75880 2440
rect 77392 2388 77444 2440
rect 78036 2388 78088 2440
rect 79508 2431 79560 2440
rect 79508 2397 79517 2431
rect 79517 2397 79551 2431
rect 79551 2397 79560 2431
rect 79508 2388 79560 2397
rect 80520 2388 80572 2440
rect 81348 2431 81400 2440
rect 81348 2397 81357 2431
rect 81357 2397 81391 2431
rect 81391 2397 81400 2431
rect 81348 2388 81400 2397
rect 86316 2456 86368 2508
rect 89536 2456 89588 2508
rect 81532 2320 81584 2372
rect 81992 2388 82044 2440
rect 83096 2388 83148 2440
rect 84568 2431 84620 2440
rect 84568 2397 84577 2431
rect 84577 2397 84611 2431
rect 84611 2397 84620 2431
rect 84568 2388 84620 2397
rect 85304 2431 85356 2440
rect 85304 2397 85313 2431
rect 85313 2397 85347 2431
rect 85347 2397 85356 2431
rect 85304 2388 85356 2397
rect 85672 2388 85724 2440
rect 87604 2388 87656 2440
rect 87696 2431 87748 2440
rect 87696 2397 87705 2431
rect 87705 2397 87739 2431
rect 87739 2397 87748 2431
rect 87696 2388 87748 2397
rect 88984 2431 89036 2440
rect 88984 2397 88993 2431
rect 88993 2397 89027 2431
rect 89027 2397 89036 2431
rect 88984 2388 89036 2397
rect 89168 2388 89220 2440
rect 90456 2431 90508 2440
rect 90456 2397 90465 2431
rect 90465 2397 90499 2431
rect 90499 2397 90508 2431
rect 90456 2388 90508 2397
rect 76840 2252 76892 2304
rect 77116 2252 77168 2304
rect 77392 2252 77444 2304
rect 77760 2295 77812 2304
rect 77760 2261 77769 2295
rect 77769 2261 77803 2295
rect 77803 2261 77812 2295
rect 77760 2252 77812 2261
rect 78588 2252 78640 2304
rect 79232 2252 79284 2304
rect 82084 2320 82136 2372
rect 91468 2388 91520 2440
rect 92112 2388 92164 2440
rect 92756 2388 92808 2440
rect 94320 2431 94372 2440
rect 94320 2397 94329 2431
rect 94329 2397 94363 2431
rect 94363 2397 94372 2431
rect 94320 2388 94372 2397
rect 92296 2320 92348 2372
rect 99656 2388 99708 2440
rect 100484 2388 100536 2440
rect 100668 2388 100720 2440
rect 104532 2388 104584 2440
rect 104900 2388 104952 2440
rect 106004 2431 106056 2440
rect 106004 2397 106013 2431
rect 106013 2397 106047 2431
rect 106047 2397 106056 2431
rect 106004 2388 106056 2397
rect 107476 2388 107528 2440
rect 94688 2320 94740 2372
rect 96620 2320 96672 2372
rect 97908 2320 97960 2372
rect 99196 2320 99248 2372
rect 101128 2320 101180 2372
rect 103060 2320 103112 2372
rect 104992 2320 105044 2372
rect 108120 2388 108172 2440
rect 108304 2431 108356 2440
rect 108304 2397 108313 2431
rect 108313 2397 108347 2431
rect 108347 2397 108356 2431
rect 108304 2388 108356 2397
rect 84016 2252 84068 2304
rect 85028 2252 85080 2304
rect 85488 2252 85540 2304
rect 88248 2252 88300 2304
rect 89168 2252 89220 2304
rect 90180 2252 90232 2304
rect 91560 2295 91612 2304
rect 91560 2261 91569 2295
rect 91569 2261 91603 2295
rect 91603 2261 91612 2295
rect 91560 2252 91612 2261
rect 92204 2295 92256 2304
rect 92204 2261 92213 2295
rect 92213 2261 92247 2295
rect 92247 2261 92256 2295
rect 92204 2252 92256 2261
rect 93032 2295 93084 2304
rect 93032 2261 93041 2295
rect 93041 2261 93075 2295
rect 93075 2261 93084 2295
rect 93032 2252 93084 2261
rect 94044 2252 94096 2304
rect 94964 2295 95016 2304
rect 94964 2261 94973 2295
rect 94973 2261 95007 2295
rect 95007 2261 95016 2295
rect 94964 2252 95016 2261
rect 95976 2252 96028 2304
rect 97080 2295 97132 2304
rect 97080 2261 97089 2295
rect 97089 2261 97123 2295
rect 97123 2261 97132 2295
rect 97080 2252 97132 2261
rect 98184 2295 98236 2304
rect 98184 2261 98193 2295
rect 98193 2261 98227 2295
rect 98227 2261 98236 2295
rect 98184 2252 98236 2261
rect 104348 2252 104400 2304
rect 105268 2295 105320 2304
rect 105268 2261 105277 2295
rect 105277 2261 105311 2295
rect 105311 2261 105320 2295
rect 105268 2252 105320 2261
rect 105636 2252 105688 2304
rect 106924 2252 106976 2304
rect 108856 2320 108908 2372
rect 110052 2456 110104 2508
rect 110788 2388 110840 2440
rect 112076 2388 112128 2440
rect 112444 2431 112496 2440
rect 112444 2397 112453 2431
rect 112453 2397 112487 2431
rect 112487 2397 112496 2431
rect 112444 2388 112496 2397
rect 113640 2431 113692 2440
rect 113640 2397 113649 2431
rect 113649 2397 113683 2431
rect 113683 2397 113692 2431
rect 113640 2388 113692 2397
rect 114008 2388 114060 2440
rect 115296 2388 115348 2440
rect 118148 2388 118200 2440
rect 116400 2363 116452 2372
rect 116400 2329 116409 2363
rect 116409 2329 116443 2363
rect 116443 2329 116452 2363
rect 116400 2320 116452 2329
rect 116584 2320 116636 2372
rect 109960 2295 110012 2304
rect 109960 2261 109969 2295
rect 109969 2261 110003 2295
rect 110003 2261 110012 2295
rect 109960 2252 110012 2261
rect 113364 2252 113416 2304
rect 115572 2295 115624 2304
rect 115572 2261 115581 2295
rect 115581 2261 115615 2295
rect 115615 2261 115624 2295
rect 115572 2252 115624 2261
rect 116492 2295 116544 2304
rect 116492 2261 116501 2295
rect 116501 2261 116535 2295
rect 116535 2261 116544 2295
rect 116492 2252 116544 2261
rect 30398 2150 30450 2202
rect 30462 2150 30514 2202
rect 30526 2150 30578 2202
rect 30590 2150 30642 2202
rect 30654 2150 30706 2202
rect 59846 2150 59898 2202
rect 59910 2150 59962 2202
rect 59974 2150 60026 2202
rect 60038 2150 60090 2202
rect 60102 2150 60154 2202
rect 89294 2150 89346 2202
rect 89358 2150 89410 2202
rect 89422 2150 89474 2202
rect 89486 2150 89538 2202
rect 89550 2150 89602 2202
rect 10140 2048 10192 2100
rect 60648 2048 60700 2100
rect 60740 2048 60792 2100
rect 66076 2048 66128 2100
rect 66812 2048 66864 2100
rect 1676 1980 1728 2032
rect 28264 1980 28316 2032
rect 28448 1980 28500 2032
rect 29828 1980 29880 2032
rect 30748 1980 30800 2032
rect 37740 1980 37792 2032
rect 38660 1980 38712 2032
rect 60924 1980 60976 2032
rect 61016 1980 61068 2032
rect 63500 1980 63552 2032
rect 67180 2048 67232 2100
rect 73528 2048 73580 2100
rect 73620 2048 73672 2100
rect 118056 2048 118108 2100
rect 116492 1980 116544 2032
rect 12532 1912 12584 1964
rect 40500 1912 40552 1964
rect 40868 1912 40920 1964
rect 7380 1844 7432 1896
rect 31392 1844 31444 1896
rect 31576 1844 31628 1896
rect 38476 1844 38528 1896
rect 46664 1912 46716 1964
rect 55220 1912 55272 1964
rect 55312 1912 55364 1964
rect 60740 1912 60792 1964
rect 60832 1912 60884 1964
rect 73896 1912 73948 1964
rect 73988 1912 74040 1964
rect 105268 1912 105320 1964
rect 70952 1844 71004 1896
rect 71044 1844 71096 1896
rect 75368 1844 75420 1896
rect 75552 1844 75604 1896
rect 77208 1844 77260 1896
rect 77392 1844 77444 1896
rect 109776 1844 109828 1896
rect 15752 1776 15804 1828
rect 42708 1776 42760 1828
rect 45928 1776 45980 1828
rect 17500 1708 17552 1760
rect 27712 1708 27764 1760
rect 29736 1708 29788 1760
rect 49700 1708 49752 1760
rect 51540 1776 51592 1828
rect 58164 1776 58216 1828
rect 58256 1776 58308 1828
rect 89536 1776 89588 1828
rect 89628 1776 89680 1828
rect 51632 1708 51684 1760
rect 51816 1708 51868 1760
rect 3516 1640 3568 1692
rect 55956 1640 56008 1692
rect 56416 1640 56468 1692
rect 58072 1640 58124 1692
rect 66904 1640 66956 1692
rect 71320 1640 71372 1692
rect 71872 1640 71924 1692
rect 73988 1640 74040 1692
rect 74080 1640 74132 1692
rect 75092 1640 75144 1692
rect 76840 1708 76892 1760
rect 91560 1708 91612 1760
rect 94780 1776 94832 1828
rect 100668 1708 100720 1760
rect 100852 1776 100904 1828
rect 106004 1776 106056 1828
rect 112444 1708 112496 1760
rect 77760 1640 77812 1692
rect 77852 1640 77904 1692
rect 98184 1640 98236 1692
rect 7196 1572 7248 1624
rect 45560 1572 45612 1624
rect 45652 1572 45704 1624
rect 52000 1572 52052 1624
rect 53104 1572 53156 1624
rect 109960 1572 110012 1624
rect 12348 1504 12400 1556
rect 18236 1436 18288 1488
rect 30748 1436 30800 1488
rect 31668 1436 31720 1488
rect 89352 1436 89404 1488
rect 89628 1504 89680 1556
rect 89720 1504 89772 1556
rect 89812 1504 89864 1556
rect 94320 1504 94372 1556
rect 97816 1504 97868 1556
rect 100852 1504 100904 1556
rect 94964 1436 95016 1488
rect 7012 1368 7064 1420
rect 80060 1368 80112 1420
rect 80152 1368 80204 1420
rect 86500 1368 86552 1420
rect 86592 1368 86644 1420
rect 89444 1368 89496 1420
rect 89536 1368 89588 1420
rect 97080 1368 97132 1420
rect 107568 1368 107620 1420
rect 108304 1368 108356 1420
rect 28908 1300 28960 1352
rect 93032 1300 93084 1352
rect 22468 1232 22520 1284
rect 31668 1232 31720 1284
rect 41788 1232 41840 1284
rect 90456 1232 90508 1284
rect 47952 1164 48004 1216
rect 81348 1164 81400 1216
rect 86500 1164 86552 1216
rect 89536 1164 89588 1216
rect 57152 1096 57204 1148
rect 87696 1096 87748 1148
<< metal2 >>
rect 18 29200 74 30000
rect 662 29322 718 30000
rect 662 29294 1072 29322
rect 662 29200 718 29294
rect 32 26246 60 29200
rect 1044 27130 1072 29294
rect 1306 29200 1362 30000
rect 2594 29322 2650 30000
rect 2424 29294 2650 29322
rect 1214 28656 1270 28665
rect 1214 28591 1270 28600
rect 1032 27124 1084 27130
rect 1032 27066 1084 27072
rect 1228 26450 1256 28591
rect 1320 26994 1348 29200
rect 2424 27538 2452 29294
rect 2594 29200 2650 29294
rect 3238 29322 3294 30000
rect 4526 29322 4582 30000
rect 5170 29322 5226 30000
rect 6458 29322 6514 30000
rect 3238 29294 3648 29322
rect 3238 29200 3294 29294
rect 2778 27976 2834 27985
rect 2778 27911 2834 27920
rect 2412 27532 2464 27538
rect 2412 27474 2464 27480
rect 2688 27464 2740 27470
rect 2688 27406 2740 27412
rect 1400 27328 1452 27334
rect 1400 27270 1452 27276
rect 1308 26988 1360 26994
rect 1308 26930 1360 26936
rect 1412 26625 1440 27270
rect 1676 26920 1728 26926
rect 1676 26862 1728 26868
rect 1398 26616 1454 26625
rect 1688 26586 1716 26862
rect 1398 26551 1454 26560
rect 1676 26580 1728 26586
rect 1676 26522 1728 26528
rect 1216 26444 1268 26450
rect 1216 26386 1268 26392
rect 20 26240 72 26246
rect 20 26182 72 26188
rect 1400 26036 1452 26042
rect 1400 25978 1452 25984
rect 1412 25945 1440 25978
rect 1398 25936 1454 25945
rect 1398 25871 1454 25880
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1412 24585 1440 24686
rect 1398 24576 1454 24585
rect 1398 24511 1454 24520
rect 2700 24206 2728 27406
rect 2792 26518 2820 27911
rect 3620 27470 3648 29294
rect 4526 29294 4660 29322
rect 4526 29200 4582 29294
rect 3608 27464 3660 27470
rect 3608 27406 3660 27412
rect 4436 27396 4488 27402
rect 4436 27338 4488 27344
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 2780 26512 2832 26518
rect 2780 26454 2832 26460
rect 2884 26246 2912 26930
rect 2964 26852 3016 26858
rect 2964 26794 3016 26800
rect 2872 26240 2924 26246
rect 2872 26182 2924 26188
rect 2976 24206 3004 26794
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1676 24200 1728 24206
rect 1676 24142 1728 24148
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 1412 23905 1440 24142
rect 1492 24064 1544 24070
rect 1492 24006 1544 24012
rect 1398 23896 1454 23905
rect 1398 23831 1454 23840
rect 1400 23520 1452 23526
rect 1400 23462 1452 23468
rect 1412 23225 1440 23462
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1400 21888 1452 21894
rect 1398 21856 1400 21865
rect 1452 21856 1454 21865
rect 1398 21791 1454 21800
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21185 1440 21490
rect 1398 21176 1454 21185
rect 1398 21111 1454 21120
rect 1398 19816 1454 19825
rect 1398 19751 1454 19760
rect 1412 19718 1440 19751
rect 1400 19712 1452 19718
rect 1400 19654 1452 19660
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 1412 18465 1440 18566
rect 1398 18456 1454 18465
rect 1398 18391 1454 18400
rect 1398 17096 1454 17105
rect 1398 17031 1400 17040
rect 1452 17031 1454 17040
rect 1400 17002 1452 17008
rect 1400 15360 1452 15366
rect 1400 15302 1452 15308
rect 1412 15065 1440 15302
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1398 14376 1454 14385
rect 1398 14311 1454 14320
rect 1412 14278 1440 14311
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1412 12345 1440 12582
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1504 11762 1532 24006
rect 1688 22982 1716 24142
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 21146 1624 21286
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1596 16425 1624 16526
rect 1582 16416 1638 16425
rect 1582 16351 1638 16360
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1398 11656 1454 11665
rect 1398 11591 1400 11600
rect 1452 11591 1454 11600
rect 1400 11562 1452 11568
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 10305 1440 10406
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 8265 1440 8298
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7585 1440 7822
rect 1398 7576 1454 7585
rect 1398 7511 1454 7520
rect 1398 6216 1454 6225
rect 1398 6151 1400 6160
rect 1452 6151 1454 6160
rect 1400 6122 1452 6128
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1412 4865 1440 5170
rect 1398 4856 1454 4865
rect 1398 4791 1454 4800
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 664 3460 716 3466
rect 664 3402 716 3408
rect 20 2916 72 2922
rect 20 2858 72 2864
rect 32 800 60 2858
rect 676 800 704 3402
rect 1308 3392 1360 3398
rect 1308 3334 1360 3340
rect 1320 800 1348 3334
rect 1412 2825 1440 4082
rect 1504 4010 1532 9998
rect 1780 4146 1808 23666
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1872 19145 1900 19314
rect 1858 19136 1914 19145
rect 1858 19071 1914 19080
rect 2228 18692 2280 18698
rect 2228 18634 2280 18640
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1964 16998 1992 17138
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1964 16454 1992 16934
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1872 13025 1900 13194
rect 1858 13016 1914 13025
rect 1858 12951 1914 12960
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1872 9625 1900 9930
rect 1858 9616 1914 9625
rect 1858 9551 1914 9560
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1964 6118 1992 6258
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1872 5545 1900 5578
rect 1858 5536 1914 5545
rect 1858 5471 1914 5480
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1964 4078 1992 6054
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1492 4004 1544 4010
rect 1492 3946 1544 3952
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 1584 3528 1636 3534
rect 1582 3496 1584 3505
rect 1636 3496 1638 3505
rect 1582 3431 1638 3440
rect 2148 3194 2176 3946
rect 2240 3534 2268 18634
rect 3528 16658 3556 26930
rect 4448 25498 4476 27338
rect 4632 27130 4660 29294
rect 5000 29294 5226 29322
rect 5000 27538 5028 29294
rect 5170 29200 5226 29294
rect 6380 29294 6514 29322
rect 6380 27538 6408 29294
rect 6458 29200 6514 29294
rect 7102 29200 7158 30000
rect 7746 29322 7802 30000
rect 7746 29294 7880 29322
rect 7746 29200 7802 29294
rect 4988 27532 5040 27538
rect 4988 27474 5040 27480
rect 6368 27532 6420 27538
rect 6368 27474 6420 27480
rect 7116 27470 7144 29200
rect 6644 27464 6696 27470
rect 6644 27406 6696 27412
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 4436 25492 4488 25498
rect 4436 25434 4488 25440
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2424 14414 2452 14962
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 6914 2452 14350
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2516 10266 2544 10610
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2608 6914 2636 16458
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2700 10062 2728 11086
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 4816 7206 4844 26930
rect 6656 26450 6684 27406
rect 7852 27130 7880 29294
rect 9034 29200 9090 30000
rect 9678 29200 9734 30000
rect 10966 29200 11022 30000
rect 11610 29200 11666 30000
rect 12254 29322 12310 30000
rect 13542 29322 13598 30000
rect 14186 29322 14242 30000
rect 12254 29294 12388 29322
rect 12254 29200 12310 29294
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 6644 26444 6696 26450
rect 6644 26386 6696 26392
rect 9048 26246 9076 29200
rect 9588 27600 9640 27606
rect 9588 27542 9640 27548
rect 9404 27396 9456 27402
rect 9404 27338 9456 27344
rect 9416 26858 9444 27338
rect 9404 26852 9456 26858
rect 9404 26794 9456 26800
rect 9600 26790 9628 27542
rect 9692 27130 9720 29200
rect 9864 27872 9916 27878
rect 9864 27814 9916 27820
rect 9876 27606 9904 27814
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 10980 27452 11008 29200
rect 11060 27464 11112 27470
rect 10980 27424 11060 27452
rect 11060 27406 11112 27412
rect 10324 27396 10376 27402
rect 10324 27338 10376 27344
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 9588 26784 9640 26790
rect 9588 26726 9640 26732
rect 9036 26240 9088 26246
rect 9036 26182 9088 26188
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 2424 6886 2544 6914
rect 2608 6886 2728 6914
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2516 3194 2544 6886
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2608 3194 2636 4082
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1412 785 1440 2382
rect 1688 2038 1716 2382
rect 1676 2032 1728 2038
rect 1676 1974 1728 1980
rect 2608 800 2636 2994
rect 2700 2446 2728 6886
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2792 1465 2820 3062
rect 2884 2446 2912 3334
rect 5460 3058 5488 3674
rect 7852 3058 7880 11834
rect 9232 11218 9260 22714
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 10244 3194 10272 26930
rect 10336 26246 10364 27338
rect 11624 27130 11652 29200
rect 12360 27452 12388 29294
rect 13542 29294 13768 29322
rect 13542 29200 13598 29294
rect 12440 27464 12492 27470
rect 12360 27424 12440 27452
rect 13740 27452 13768 29294
rect 14186 29294 14320 29322
rect 14186 29200 14242 29294
rect 13820 27464 13872 27470
rect 13740 27424 13820 27452
rect 12440 27406 12492 27412
rect 13820 27406 13872 27412
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 12532 27328 12584 27334
rect 12532 27270 12584 27276
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11992 27062 12020 27270
rect 11980 27056 12032 27062
rect 11980 26998 12032 27004
rect 10508 26852 10560 26858
rect 10508 26794 10560 26800
rect 10324 26240 10376 26246
rect 10324 26182 10376 26188
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15162 10456 15438
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10520 6914 10548 26794
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10888 15026 10916 15302
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10428 6886 10548 6914
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3252 800 3280 2382
rect 3528 1698 3556 2994
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 3516 1692 3568 1698
rect 3516 1634 3568 1640
rect 4540 800 4568 2382
rect 5184 800 5212 2790
rect 5828 800 5856 2790
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7024 1426 7052 2246
rect 7012 1420 7064 1426
rect 7012 1362 7064 1368
rect 7116 800 7144 2790
rect 7208 1630 7236 2994
rect 7392 1902 7420 2994
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7380 1896 7432 1902
rect 7380 1838 7432 1844
rect 7196 1624 7248 1630
rect 7196 1566 7248 1572
rect 7760 800 7788 2926
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9048 800 9076 2382
rect 9692 800 9720 2518
rect 10428 2446 10456 6886
rect 10888 2650 10916 14962
rect 11716 12306 11744 22918
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10152 2106 10180 2246
rect 10140 2100 10192 2106
rect 10140 2042 10192 2048
rect 10980 800 11008 2314
rect 11624 800 11652 2382
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 800 12296 2246
rect 12360 1562 12388 2994
rect 12544 1970 12572 27270
rect 14292 26994 14320 29294
rect 15474 29200 15530 30000
rect 16118 29200 16174 30000
rect 17406 29322 17462 30000
rect 17236 29294 17462 29322
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 14462 27296 14518 27305
rect 14462 27231 14518 27240
rect 14476 27062 14504 27231
rect 14464 27056 14516 27062
rect 15212 27033 15240 27338
rect 15488 27062 15516 29200
rect 15674 27772 15982 27781
rect 15674 27770 15680 27772
rect 15736 27770 15760 27772
rect 15816 27770 15840 27772
rect 15896 27770 15920 27772
rect 15976 27770 15982 27772
rect 15736 27718 15738 27770
rect 15918 27718 15920 27770
rect 15674 27716 15680 27718
rect 15736 27716 15760 27718
rect 15816 27716 15840 27718
rect 15896 27716 15920 27718
rect 15976 27716 15982 27718
rect 15674 27707 15982 27716
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 15476 27056 15528 27062
rect 14464 26998 14516 27004
rect 15198 27024 15254 27033
rect 14280 26988 14332 26994
rect 15476 26998 15528 27004
rect 16040 27010 16068 27406
rect 16132 27402 16160 29200
rect 17132 27872 17184 27878
rect 17132 27814 17184 27820
rect 17144 27674 17172 27814
rect 17132 27668 17184 27674
rect 17132 27610 17184 27616
rect 17040 27600 17092 27606
rect 17040 27542 17092 27548
rect 16120 27396 16172 27402
rect 16120 27338 16172 27344
rect 16212 27396 16264 27402
rect 16212 27338 16264 27344
rect 16224 27305 16252 27338
rect 16210 27296 16266 27305
rect 16210 27231 16266 27240
rect 16040 26982 16160 27010
rect 15198 26959 15254 26968
rect 14280 26930 14332 26936
rect 16028 26852 16080 26858
rect 16028 26794 16080 26800
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15580 26518 15608 26726
rect 15674 26684 15982 26693
rect 15674 26682 15680 26684
rect 15736 26682 15760 26684
rect 15816 26682 15840 26684
rect 15896 26682 15920 26684
rect 15976 26682 15982 26684
rect 15736 26630 15738 26682
rect 15918 26630 15920 26682
rect 15674 26628 15680 26630
rect 15736 26628 15760 26630
rect 15816 26628 15840 26630
rect 15896 26628 15920 26630
rect 15976 26628 15982 26630
rect 15674 26619 15982 26628
rect 15568 26512 15620 26518
rect 15568 26454 15620 26460
rect 15674 25596 15982 25605
rect 15674 25594 15680 25596
rect 15736 25594 15760 25596
rect 15816 25594 15840 25596
rect 15896 25594 15920 25596
rect 15976 25594 15982 25596
rect 15736 25542 15738 25594
rect 15918 25542 15920 25594
rect 15674 25540 15680 25542
rect 15736 25540 15760 25542
rect 15816 25540 15840 25542
rect 15896 25540 15920 25542
rect 15976 25540 15982 25542
rect 15674 25531 15982 25540
rect 15674 24508 15982 24517
rect 15674 24506 15680 24508
rect 15736 24506 15760 24508
rect 15816 24506 15840 24508
rect 15896 24506 15920 24508
rect 15976 24506 15982 24508
rect 15736 24454 15738 24506
rect 15918 24454 15920 24506
rect 15674 24452 15680 24454
rect 15736 24452 15760 24454
rect 15816 24452 15840 24454
rect 15896 24452 15920 24454
rect 15976 24452 15982 24454
rect 15674 24443 15982 24452
rect 15674 23420 15982 23429
rect 15674 23418 15680 23420
rect 15736 23418 15760 23420
rect 15816 23418 15840 23420
rect 15896 23418 15920 23420
rect 15976 23418 15982 23420
rect 15736 23366 15738 23418
rect 15918 23366 15920 23418
rect 15674 23364 15680 23366
rect 15736 23364 15760 23366
rect 15816 23364 15840 23366
rect 15896 23364 15920 23366
rect 15976 23364 15982 23366
rect 15674 23355 15982 23364
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12636 2446 12664 2790
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 12532 1964 12584 1970
rect 12532 1906 12584 1912
rect 12348 1556 12400 1562
rect 12348 1498 12400 1504
rect 13556 800 13584 2314
rect 14200 800 14228 2994
rect 14660 2650 14688 22918
rect 15674 22332 15982 22341
rect 15674 22330 15680 22332
rect 15736 22330 15760 22332
rect 15816 22330 15840 22332
rect 15896 22330 15920 22332
rect 15976 22330 15982 22332
rect 15736 22278 15738 22330
rect 15918 22278 15920 22330
rect 15674 22276 15680 22278
rect 15736 22276 15760 22278
rect 15816 22276 15840 22278
rect 15896 22276 15920 22278
rect 15976 22276 15982 22278
rect 15674 22267 15982 22276
rect 15674 21244 15982 21253
rect 15674 21242 15680 21244
rect 15736 21242 15760 21244
rect 15816 21242 15840 21244
rect 15896 21242 15920 21244
rect 15976 21242 15982 21244
rect 15736 21190 15738 21242
rect 15918 21190 15920 21242
rect 15674 21188 15680 21190
rect 15736 21188 15760 21190
rect 15816 21188 15840 21190
rect 15896 21188 15920 21190
rect 15976 21188 15982 21190
rect 15674 21179 15982 21188
rect 15674 20156 15982 20165
rect 15674 20154 15680 20156
rect 15736 20154 15760 20156
rect 15816 20154 15840 20156
rect 15896 20154 15920 20156
rect 15976 20154 15982 20156
rect 15736 20102 15738 20154
rect 15918 20102 15920 20154
rect 15674 20100 15680 20102
rect 15736 20100 15760 20102
rect 15816 20100 15840 20102
rect 15896 20100 15920 20102
rect 15976 20100 15982 20102
rect 15674 20091 15982 20100
rect 15674 19068 15982 19077
rect 15674 19066 15680 19068
rect 15736 19066 15760 19068
rect 15816 19066 15840 19068
rect 15896 19066 15920 19068
rect 15976 19066 15982 19068
rect 15736 19014 15738 19066
rect 15918 19014 15920 19066
rect 15674 19012 15680 19014
rect 15736 19012 15760 19014
rect 15816 19012 15840 19014
rect 15896 19012 15920 19014
rect 15976 19012 15982 19014
rect 15674 19003 15982 19012
rect 15674 17980 15982 17989
rect 15674 17978 15680 17980
rect 15736 17978 15760 17980
rect 15816 17978 15840 17980
rect 15896 17978 15920 17980
rect 15976 17978 15982 17980
rect 15736 17926 15738 17978
rect 15918 17926 15920 17978
rect 15674 17924 15680 17926
rect 15736 17924 15760 17926
rect 15816 17924 15840 17926
rect 15896 17924 15920 17926
rect 15976 17924 15982 17926
rect 15674 17915 15982 17924
rect 15674 16892 15982 16901
rect 15674 16890 15680 16892
rect 15736 16890 15760 16892
rect 15816 16890 15840 16892
rect 15896 16890 15920 16892
rect 15976 16890 15982 16892
rect 15736 16838 15738 16890
rect 15918 16838 15920 16890
rect 15674 16836 15680 16838
rect 15736 16836 15760 16838
rect 15816 16836 15840 16838
rect 15896 16836 15920 16838
rect 15976 16836 15982 16838
rect 15674 16827 15982 16836
rect 15674 15804 15982 15813
rect 15674 15802 15680 15804
rect 15736 15802 15760 15804
rect 15816 15802 15840 15804
rect 15896 15802 15920 15804
rect 15976 15802 15982 15804
rect 15736 15750 15738 15802
rect 15918 15750 15920 15802
rect 15674 15748 15680 15750
rect 15736 15748 15760 15750
rect 15816 15748 15840 15750
rect 15896 15748 15920 15750
rect 15976 15748 15982 15750
rect 15674 15739 15982 15748
rect 15674 14716 15982 14725
rect 15674 14714 15680 14716
rect 15736 14714 15760 14716
rect 15816 14714 15840 14716
rect 15896 14714 15920 14716
rect 15976 14714 15982 14716
rect 15736 14662 15738 14714
rect 15918 14662 15920 14714
rect 15674 14660 15680 14662
rect 15736 14660 15760 14662
rect 15816 14660 15840 14662
rect 15896 14660 15920 14662
rect 15976 14660 15982 14662
rect 15674 14651 15982 14660
rect 15674 13628 15982 13637
rect 15674 13626 15680 13628
rect 15736 13626 15760 13628
rect 15816 13626 15840 13628
rect 15896 13626 15920 13628
rect 15976 13626 15982 13628
rect 15736 13574 15738 13626
rect 15918 13574 15920 13626
rect 15674 13572 15680 13574
rect 15736 13572 15760 13574
rect 15816 13572 15840 13574
rect 15896 13572 15920 13574
rect 15976 13572 15982 13574
rect 15674 13563 15982 13572
rect 16040 13258 16068 26794
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 15674 12540 15982 12549
rect 15674 12538 15680 12540
rect 15736 12538 15760 12540
rect 15816 12538 15840 12540
rect 15896 12538 15920 12540
rect 15976 12538 15982 12540
rect 15736 12486 15738 12538
rect 15918 12486 15920 12538
rect 15674 12484 15680 12486
rect 15736 12484 15760 12486
rect 15816 12484 15840 12486
rect 15896 12484 15920 12486
rect 15976 12484 15982 12486
rect 15674 12475 15982 12484
rect 15674 11452 15982 11461
rect 15674 11450 15680 11452
rect 15736 11450 15760 11452
rect 15816 11450 15840 11452
rect 15896 11450 15920 11452
rect 15976 11450 15982 11452
rect 15736 11398 15738 11450
rect 15918 11398 15920 11450
rect 15674 11396 15680 11398
rect 15736 11396 15760 11398
rect 15816 11396 15840 11398
rect 15896 11396 15920 11398
rect 15976 11396 15982 11398
rect 15674 11387 15982 11396
rect 15674 10364 15982 10373
rect 15674 10362 15680 10364
rect 15736 10362 15760 10364
rect 15816 10362 15840 10364
rect 15896 10362 15920 10364
rect 15976 10362 15982 10364
rect 15736 10310 15738 10362
rect 15918 10310 15920 10362
rect 15674 10308 15680 10310
rect 15736 10308 15760 10310
rect 15816 10308 15840 10310
rect 15896 10308 15920 10310
rect 15976 10308 15982 10310
rect 15674 10299 15982 10308
rect 15674 9276 15982 9285
rect 15674 9274 15680 9276
rect 15736 9274 15760 9276
rect 15816 9274 15840 9276
rect 15896 9274 15920 9276
rect 15976 9274 15982 9276
rect 15736 9222 15738 9274
rect 15918 9222 15920 9274
rect 15674 9220 15680 9222
rect 15736 9220 15760 9222
rect 15816 9220 15840 9222
rect 15896 9220 15920 9222
rect 15976 9220 15982 9222
rect 15674 9211 15982 9220
rect 15674 8188 15982 8197
rect 15674 8186 15680 8188
rect 15736 8186 15760 8188
rect 15816 8186 15840 8188
rect 15896 8186 15920 8188
rect 15976 8186 15982 8188
rect 15736 8134 15738 8186
rect 15918 8134 15920 8186
rect 15674 8132 15680 8134
rect 15736 8132 15760 8134
rect 15816 8132 15840 8134
rect 15896 8132 15920 8134
rect 15976 8132 15982 8134
rect 15674 8123 15982 8132
rect 15674 7100 15982 7109
rect 15674 7098 15680 7100
rect 15736 7098 15760 7100
rect 15816 7098 15840 7100
rect 15896 7098 15920 7100
rect 15976 7098 15982 7100
rect 15736 7046 15738 7098
rect 15918 7046 15920 7098
rect 15674 7044 15680 7046
rect 15736 7044 15760 7046
rect 15816 7044 15840 7046
rect 15896 7044 15920 7046
rect 15976 7044 15982 7046
rect 15674 7035 15982 7044
rect 15674 6012 15982 6021
rect 15674 6010 15680 6012
rect 15736 6010 15760 6012
rect 15816 6010 15840 6012
rect 15896 6010 15920 6012
rect 15976 6010 15982 6012
rect 15736 5958 15738 6010
rect 15918 5958 15920 6010
rect 15674 5956 15680 5958
rect 15736 5956 15760 5958
rect 15816 5956 15840 5958
rect 15896 5956 15920 5958
rect 15976 5956 15982 5958
rect 15674 5947 15982 5956
rect 15674 4924 15982 4933
rect 15674 4922 15680 4924
rect 15736 4922 15760 4924
rect 15816 4922 15840 4924
rect 15896 4922 15920 4924
rect 15976 4922 15982 4924
rect 15736 4870 15738 4922
rect 15918 4870 15920 4922
rect 15674 4868 15680 4870
rect 15736 4868 15760 4870
rect 15816 4868 15840 4870
rect 15896 4868 15920 4870
rect 15976 4868 15982 4870
rect 15674 4859 15982 4868
rect 15674 3836 15982 3845
rect 15674 3834 15680 3836
rect 15736 3834 15760 3836
rect 15816 3834 15840 3836
rect 15896 3834 15920 3836
rect 15976 3834 15982 3836
rect 15736 3782 15738 3834
rect 15918 3782 15920 3834
rect 15674 3780 15680 3782
rect 15736 3780 15760 3782
rect 15816 3780 15840 3782
rect 15896 3780 15920 3782
rect 15976 3780 15982 3782
rect 15674 3771 15982 3780
rect 15674 2748 15982 2757
rect 15674 2746 15680 2748
rect 15736 2746 15760 2748
rect 15816 2746 15840 2748
rect 15896 2746 15920 2748
rect 15976 2746 15982 2748
rect 15736 2694 15738 2746
rect 15918 2694 15920 2746
rect 15674 2692 15680 2694
rect 15736 2692 15760 2694
rect 15816 2692 15840 2694
rect 15896 2692 15920 2694
rect 15976 2692 15982 2694
rect 15674 2683 15982 2692
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 16132 2514 16160 26982
rect 17052 26858 17080 27542
rect 17236 27470 17264 29294
rect 17406 29200 17462 29294
rect 18050 29200 18106 30000
rect 18694 29200 18750 30000
rect 19982 29322 20038 30000
rect 19982 29294 20208 29322
rect 19982 29200 20038 29294
rect 18064 27470 18092 29200
rect 18708 27606 18736 29200
rect 19800 27872 19852 27878
rect 19800 27814 19852 27820
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 17224 27464 17276 27470
rect 17224 27406 17276 27412
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 19352 27402 19380 27542
rect 19340 27396 19392 27402
rect 19340 27338 19392 27344
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17316 27328 17368 27334
rect 17316 27270 17368 27276
rect 17144 27062 17172 27270
rect 17132 27056 17184 27062
rect 17132 26998 17184 27004
rect 17040 26852 17092 26858
rect 17040 26794 17092 26800
rect 16854 2544 16910 2553
rect 16120 2508 16172 2514
rect 16854 2479 16910 2488
rect 16120 2450 16172 2456
rect 16868 2446 16896 2479
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15488 800 15516 2246
rect 15764 1834 15792 2382
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 15752 1828 15804 1834
rect 15752 1770 15804 1776
rect 16132 800 16160 2246
rect 17328 1601 17356 27270
rect 19708 27056 19760 27062
rect 19708 26998 19760 27004
rect 19720 26761 19748 26998
rect 19812 26994 19840 27814
rect 20180 27470 20208 29294
rect 20626 29200 20682 30000
rect 21914 29322 21970 30000
rect 22558 29322 22614 30000
rect 21914 29294 22048 29322
rect 21914 29200 21970 29294
rect 20168 27464 20220 27470
rect 20168 27406 20220 27412
rect 20352 27464 20404 27470
rect 20352 27406 20404 27412
rect 20536 27464 20588 27470
rect 20640 27452 20668 29200
rect 21178 27704 21234 27713
rect 21178 27639 21234 27648
rect 21088 27464 21140 27470
rect 20640 27424 20852 27452
rect 20536 27406 20588 27412
rect 19800 26988 19852 26994
rect 19800 26930 19852 26936
rect 19706 26752 19762 26761
rect 19706 26687 19762 26696
rect 20364 26489 20392 27406
rect 20548 26858 20576 27406
rect 20824 27334 20852 27424
rect 21088 27406 21140 27412
rect 20628 27328 20680 27334
rect 20626 27296 20628 27305
rect 20812 27328 20864 27334
rect 20680 27296 20682 27305
rect 20812 27270 20864 27276
rect 20626 27231 20682 27240
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20732 26897 20760 26930
rect 20718 26888 20774 26897
rect 20536 26852 20588 26858
rect 20718 26823 20774 26832
rect 20536 26794 20588 26800
rect 21100 26790 21128 27406
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 21192 26518 21220 27639
rect 22020 27452 22048 29294
rect 22558 29294 22692 29322
rect 22558 29200 22614 29294
rect 22664 27606 22692 29294
rect 23846 29200 23902 30000
rect 24490 29322 24546 30000
rect 24412 29294 24546 29322
rect 22652 27600 22704 27606
rect 22652 27542 22704 27548
rect 23662 27568 23718 27577
rect 22376 27532 22428 27538
rect 22376 27474 22428 27480
rect 23388 27532 23440 27538
rect 23572 27532 23624 27538
rect 23440 27492 23572 27520
rect 23388 27474 23440 27480
rect 23662 27503 23718 27512
rect 23572 27474 23624 27480
rect 22100 27464 22152 27470
rect 22020 27424 22100 27452
rect 22100 27406 22152 27412
rect 21916 27396 21968 27402
rect 21916 27338 21968 27344
rect 21928 27169 21956 27338
rect 22008 27328 22060 27334
rect 22008 27270 22060 27276
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 21914 27160 21970 27169
rect 21914 27095 21970 27104
rect 21914 27024 21970 27033
rect 21914 26959 21970 26968
rect 21928 26790 21956 26959
rect 22020 26858 22048 27270
rect 22296 27010 22324 27270
rect 22388 27062 22416 27474
rect 23676 27470 23704 27503
rect 23860 27470 23888 29200
rect 23664 27464 23716 27470
rect 23570 27432 23626 27441
rect 23664 27406 23716 27412
rect 23848 27464 23900 27470
rect 23848 27406 23900 27412
rect 23570 27367 23626 27376
rect 23584 27334 23612 27367
rect 24412 27334 24440 29294
rect 24490 29200 24546 29294
rect 25134 29322 25190 30000
rect 25134 29294 25360 29322
rect 25134 29200 25190 29294
rect 25332 27470 25360 29294
rect 26422 29200 26478 30000
rect 27066 29322 27122 30000
rect 28354 29322 28410 30000
rect 27066 29294 27384 29322
rect 27066 29200 27122 29294
rect 26436 27470 26464 29200
rect 26700 28008 26752 28014
rect 26700 27950 26752 27956
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 25148 27169 25176 27406
rect 26712 27334 26740 27950
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 26884 27396 26936 27402
rect 26884 27338 26936 27344
rect 26700 27328 26752 27334
rect 26700 27270 26752 27276
rect 25134 27160 25190 27169
rect 25134 27095 25190 27104
rect 22204 26982 22324 27010
rect 22376 27056 22428 27062
rect 26792 27056 26844 27062
rect 22376 26998 22428 27004
rect 22466 27024 22522 27033
rect 22204 26858 22232 26982
rect 22466 26959 22522 26968
rect 26790 27024 26792 27033
rect 26844 27024 26846 27033
rect 26790 26959 26846 26968
rect 22008 26852 22060 26858
rect 22008 26794 22060 26800
rect 22192 26852 22244 26858
rect 22192 26794 22244 26800
rect 22284 26852 22336 26858
rect 22284 26794 22336 26800
rect 21916 26784 21968 26790
rect 22296 26738 22324 26794
rect 21916 26726 21968 26732
rect 22112 26710 22324 26738
rect 22374 26752 22430 26761
rect 22112 26586 22140 26710
rect 22374 26687 22430 26696
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22388 26518 22416 26687
rect 22480 26625 22508 26959
rect 24124 26920 24176 26926
rect 24124 26862 24176 26868
rect 24136 26761 24164 26862
rect 26792 26852 26844 26858
rect 26792 26794 26844 26800
rect 24122 26752 24178 26761
rect 24122 26687 24178 26696
rect 22466 26616 22522 26625
rect 22466 26551 22522 26560
rect 24124 26580 24176 26586
rect 24124 26522 24176 26528
rect 21180 26512 21232 26518
rect 20350 26480 20406 26489
rect 21180 26454 21232 26460
rect 22376 26512 22428 26518
rect 22376 26454 22428 26460
rect 24136 26450 24164 26522
rect 20350 26415 20406 26424
rect 24124 26444 24176 26450
rect 24124 26386 24176 26392
rect 22376 26376 22428 26382
rect 22374 26344 22376 26353
rect 22428 26344 22430 26353
rect 22374 26279 22430 26288
rect 24490 26344 24546 26353
rect 24490 26279 24492 26288
rect 24544 26279 24546 26288
rect 24492 26250 24544 26256
rect 26804 26246 26832 26794
rect 26792 26240 26844 26246
rect 26792 26182 26844 26188
rect 26896 17678 26924 27338
rect 26976 27328 27028 27334
rect 26976 27270 27028 27276
rect 26988 27130 27016 27270
rect 26976 27124 27028 27130
rect 26976 27066 27028 27072
rect 27080 27062 27108 27814
rect 27160 27600 27212 27606
rect 27160 27542 27212 27548
rect 27068 27056 27120 27062
rect 27068 26998 27120 27004
rect 27172 26926 27200 27542
rect 27356 26994 27384 29294
rect 28092 29294 28410 29322
rect 28092 27470 28120 29294
rect 28354 29200 28410 29294
rect 28998 29200 29054 30000
rect 29642 29322 29698 30000
rect 29642 29294 29776 29322
rect 29642 29200 29698 29294
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 28908 27464 28960 27470
rect 29012 27452 29040 29200
rect 29274 27840 29330 27849
rect 29274 27775 29330 27784
rect 28960 27424 29040 27452
rect 28908 27406 28960 27412
rect 27528 27396 27580 27402
rect 27528 27338 27580 27344
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27540 26926 27568 27338
rect 29184 27124 29236 27130
rect 29184 27066 29236 27072
rect 27160 26920 27212 26926
rect 27160 26862 27212 26868
rect 27528 26920 27580 26926
rect 27528 26862 27580 26868
rect 29000 26920 29052 26926
rect 29196 26908 29224 27066
rect 29288 27062 29316 27775
rect 29552 27328 29604 27334
rect 29552 27270 29604 27276
rect 29276 27056 29328 27062
rect 29276 26998 29328 27004
rect 29564 26994 29592 27270
rect 29552 26988 29604 26994
rect 29552 26930 29604 26936
rect 29368 26920 29420 26926
rect 29196 26880 29368 26908
rect 29000 26862 29052 26868
rect 29368 26862 29420 26868
rect 27252 26852 27304 26858
rect 27252 26794 27304 26800
rect 27068 26784 27120 26790
rect 27160 26784 27212 26790
rect 27068 26726 27120 26732
rect 27158 26752 27160 26761
rect 27212 26752 27214 26761
rect 27080 26602 27108 26726
rect 27158 26687 27214 26696
rect 27264 26602 27292 26794
rect 27080 26574 27292 26602
rect 29012 26489 29040 26862
rect 29092 26852 29144 26858
rect 29552 26852 29604 26858
rect 29092 26794 29144 26800
rect 29472 26812 29552 26840
rect 28170 26480 28226 26489
rect 28170 26415 28172 26424
rect 28224 26415 28226 26424
rect 28998 26480 29054 26489
rect 28998 26415 29054 26424
rect 28172 26386 28224 26392
rect 29104 26042 29132 26794
rect 29276 26784 29328 26790
rect 29274 26752 29276 26761
rect 29328 26752 29330 26761
rect 29274 26687 29330 26696
rect 29472 26382 29500 26812
rect 29552 26794 29604 26800
rect 29748 26586 29776 29294
rect 30930 29200 30986 30000
rect 31574 29322 31630 30000
rect 31574 29294 31708 29322
rect 31574 29200 31630 29294
rect 30656 27532 30708 27538
rect 30656 27474 30708 27480
rect 30748 27532 30800 27538
rect 30748 27474 30800 27480
rect 30668 27441 30696 27474
rect 30470 27432 30526 27441
rect 30288 27396 30340 27402
rect 30470 27367 30526 27376
rect 30654 27432 30710 27441
rect 30654 27367 30710 27376
rect 30288 27338 30340 27344
rect 30102 27296 30158 27305
rect 30102 27231 30158 27240
rect 30116 26790 30144 27231
rect 30194 27160 30250 27169
rect 30194 27095 30250 27104
rect 30104 26784 30156 26790
rect 30104 26726 30156 26732
rect 29552 26580 29604 26586
rect 29552 26522 29604 26528
rect 29736 26580 29788 26586
rect 29736 26522 29788 26528
rect 29460 26376 29512 26382
rect 29460 26318 29512 26324
rect 29092 26036 29144 26042
rect 29092 25978 29144 25984
rect 29564 24954 29592 26522
rect 30208 26518 30236 27095
rect 30300 27010 30328 27338
rect 30484 27334 30512 27367
rect 30472 27328 30524 27334
rect 30472 27270 30524 27276
rect 30398 27228 30706 27237
rect 30398 27226 30404 27228
rect 30460 27226 30484 27228
rect 30540 27226 30564 27228
rect 30620 27226 30644 27228
rect 30700 27226 30706 27228
rect 30460 27174 30462 27226
rect 30642 27174 30644 27226
rect 30398 27172 30404 27174
rect 30460 27172 30484 27174
rect 30540 27172 30564 27174
rect 30620 27172 30644 27174
rect 30700 27172 30706 27174
rect 30398 27163 30706 27172
rect 30472 27124 30524 27130
rect 30472 27066 30524 27072
rect 30484 27010 30512 27066
rect 30300 26982 30512 27010
rect 30760 26994 30788 27474
rect 30944 27470 30972 29200
rect 31392 27600 31444 27606
rect 31114 27568 31170 27577
rect 31114 27503 31116 27512
rect 31168 27503 31170 27512
rect 31390 27568 31392 27577
rect 31444 27568 31446 27577
rect 31390 27503 31446 27512
rect 31116 27474 31168 27480
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 30932 27464 30984 27470
rect 30932 27406 30984 27412
rect 31680 27418 31708 29294
rect 32862 29200 32918 30000
rect 33506 29322 33562 30000
rect 34794 29322 34850 30000
rect 33336 29294 33562 29322
rect 31760 27872 31812 27878
rect 31760 27814 31812 27820
rect 32680 27872 32732 27878
rect 32680 27814 32732 27820
rect 31772 27606 31800 27814
rect 31760 27600 31812 27606
rect 31760 27542 31812 27548
rect 31864 27538 32076 27554
rect 31852 27532 32088 27538
rect 31904 27526 32036 27532
rect 31852 27474 31904 27480
rect 32036 27474 32088 27480
rect 32126 27432 32182 27441
rect 30748 26988 30800 26994
rect 30748 26930 30800 26936
rect 30104 26512 30156 26518
rect 30104 26454 30156 26460
rect 30196 26512 30248 26518
rect 30196 26454 30248 26460
rect 29644 26376 29696 26382
rect 29644 26318 29696 26324
rect 29552 24948 29604 24954
rect 29552 24890 29604 24896
rect 28816 24064 28868 24070
rect 28816 24006 28868 24012
rect 26884 17672 26936 17678
rect 26884 17614 26936 17620
rect 25412 16720 25464 16726
rect 25412 16662 25464 16668
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20640 12442 20668 12786
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 23296 12164 23348 12170
rect 23296 12106 23348 12112
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20732 3194 20760 3538
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19444 2446 19472 2586
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 19432 2440 19484 2446
rect 19984 2440 20036 2446
rect 19432 2382 19484 2388
rect 19706 2408 19762 2417
rect 17314 1592 17370 1601
rect 17314 1527 17370 1536
rect 17420 800 17448 2382
rect 18236 2372 18288 2378
rect 19984 2382 20036 2388
rect 19706 2343 19708 2352
rect 18236 2314 18288 2320
rect 19760 2343 19762 2352
rect 19708 2314 19760 2320
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 17512 1766 17540 2246
rect 17500 1760 17552 1766
rect 17500 1702 17552 1708
rect 18064 800 18092 2246
rect 18248 1494 18276 2314
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18236 1488 18288 1494
rect 18236 1430 18288 1436
rect 18708 800 18736 2246
rect 19996 800 20024 2382
rect 20640 800 20668 2994
rect 23124 2650 23152 2994
rect 23308 2650 23336 12106
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24504 3058 24532 3130
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 21928 800 21956 2382
rect 22480 1290 22508 2586
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 24676 2440 24728 2446
rect 24780 2428 24808 2790
rect 25424 2650 25452 16662
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 24860 2440 24912 2446
rect 24780 2400 24860 2428
rect 24676 2382 24728 2388
rect 24860 2382 24912 2388
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 22468 1284 22520 1290
rect 22468 1226 22520 1232
rect 22572 800 22600 2382
rect 23216 800 23244 2382
rect 24688 2310 24716 2382
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24676 2304 24728 2310
rect 24676 2246 24728 2252
rect 24504 800 24532 2246
rect 25148 800 25176 2382
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 26160 1737 26188 2246
rect 26146 1728 26202 1737
rect 26146 1663 26202 1672
rect 26436 800 26464 2790
rect 27540 2514 27568 7890
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 27632 2650 27660 2994
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 27528 2508 27580 2514
rect 27528 2450 27580 2456
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 28170 2408 28226 2417
rect 27080 800 27108 2382
rect 27160 2304 27212 2310
rect 27344 2304 27396 2310
rect 27212 2264 27344 2292
rect 27160 2246 27212 2252
rect 27344 2246 27396 2252
rect 27724 1766 27752 2382
rect 28170 2343 28226 2352
rect 28264 2372 28316 2378
rect 28184 2310 28212 2343
rect 28264 2314 28316 2320
rect 28172 2304 28224 2310
rect 28172 2246 28224 2252
rect 28276 2038 28304 2314
rect 28264 2032 28316 2038
rect 28264 1974 28316 1980
rect 27712 1760 27764 1766
rect 27712 1702 27764 1708
rect 28368 800 28396 2790
rect 28828 2650 28856 24006
rect 28908 21412 28960 21418
rect 28908 21354 28960 21360
rect 28920 3194 28948 21354
rect 29460 8424 29512 8430
rect 29460 8366 29512 8372
rect 29472 8090 29500 8366
rect 29460 8084 29512 8090
rect 29460 8026 29512 8032
rect 29656 3194 29684 26318
rect 30116 26314 30144 26454
rect 30104 26308 30156 26314
rect 30104 26250 30156 26256
rect 30398 26140 30706 26149
rect 30398 26138 30404 26140
rect 30460 26138 30484 26140
rect 30540 26138 30564 26140
rect 30620 26138 30644 26140
rect 30700 26138 30706 26140
rect 30460 26086 30462 26138
rect 30642 26086 30644 26138
rect 30398 26084 30404 26086
rect 30460 26084 30484 26086
rect 30540 26084 30564 26086
rect 30620 26084 30644 26086
rect 30700 26084 30706 26086
rect 30398 26075 30706 26084
rect 30398 25052 30706 25061
rect 30398 25050 30404 25052
rect 30460 25050 30484 25052
rect 30540 25050 30564 25052
rect 30620 25050 30644 25052
rect 30700 25050 30706 25052
rect 30460 24998 30462 25050
rect 30642 24998 30644 25050
rect 30398 24996 30404 24998
rect 30460 24996 30484 24998
rect 30540 24996 30564 24998
rect 30620 24996 30644 24998
rect 30700 24996 30706 24998
rect 30398 24987 30706 24996
rect 30398 23964 30706 23973
rect 30398 23962 30404 23964
rect 30460 23962 30484 23964
rect 30540 23962 30564 23964
rect 30620 23962 30644 23964
rect 30700 23962 30706 23964
rect 30460 23910 30462 23962
rect 30642 23910 30644 23962
rect 30398 23908 30404 23910
rect 30460 23908 30484 23910
rect 30540 23908 30564 23910
rect 30620 23908 30644 23910
rect 30700 23908 30706 23910
rect 30398 23899 30706 23908
rect 30398 22876 30706 22885
rect 30398 22874 30404 22876
rect 30460 22874 30484 22876
rect 30540 22874 30564 22876
rect 30620 22874 30644 22876
rect 30700 22874 30706 22876
rect 30460 22822 30462 22874
rect 30642 22822 30644 22874
rect 30398 22820 30404 22822
rect 30460 22820 30484 22822
rect 30540 22820 30564 22822
rect 30620 22820 30644 22822
rect 30700 22820 30706 22822
rect 30398 22811 30706 22820
rect 30852 22094 30880 27406
rect 31680 27402 32076 27418
rect 31576 27396 31628 27402
rect 31680 27396 32088 27402
rect 31680 27390 32036 27396
rect 31576 27338 31628 27344
rect 32126 27367 32128 27376
rect 32036 27338 32088 27344
rect 32180 27367 32182 27376
rect 32128 27338 32180 27344
rect 31484 27328 31536 27334
rect 31484 27270 31536 27276
rect 31496 26738 31524 27270
rect 31588 27033 31616 27338
rect 32692 27130 32720 27814
rect 32772 27396 32824 27402
rect 32772 27338 32824 27344
rect 32680 27124 32732 27130
rect 32680 27066 32732 27072
rect 31852 27056 31904 27062
rect 31574 27024 31630 27033
rect 31852 26998 31904 27004
rect 31574 26959 31630 26968
rect 31864 26874 31892 26998
rect 32036 26988 32088 26994
rect 32036 26930 32088 26936
rect 32128 26988 32180 26994
rect 32128 26930 32180 26936
rect 31404 26710 31524 26738
rect 31772 26846 31892 26874
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 31300 24744 31352 24750
rect 31300 24686 31352 24692
rect 30852 22066 30972 22094
rect 30398 21788 30706 21797
rect 30398 21786 30404 21788
rect 30460 21786 30484 21788
rect 30540 21786 30564 21788
rect 30620 21786 30644 21788
rect 30700 21786 30706 21788
rect 30460 21734 30462 21786
rect 30642 21734 30644 21786
rect 30398 21732 30404 21734
rect 30460 21732 30484 21734
rect 30540 21732 30564 21734
rect 30620 21732 30644 21734
rect 30700 21732 30706 21734
rect 30398 21723 30706 21732
rect 30398 20700 30706 20709
rect 30398 20698 30404 20700
rect 30460 20698 30484 20700
rect 30540 20698 30564 20700
rect 30620 20698 30644 20700
rect 30700 20698 30706 20700
rect 30460 20646 30462 20698
rect 30642 20646 30644 20698
rect 30398 20644 30404 20646
rect 30460 20644 30484 20646
rect 30540 20644 30564 20646
rect 30620 20644 30644 20646
rect 30700 20644 30706 20646
rect 30398 20635 30706 20644
rect 30398 19612 30706 19621
rect 30398 19610 30404 19612
rect 30460 19610 30484 19612
rect 30540 19610 30564 19612
rect 30620 19610 30644 19612
rect 30700 19610 30706 19612
rect 30460 19558 30462 19610
rect 30642 19558 30644 19610
rect 30398 19556 30404 19558
rect 30460 19556 30484 19558
rect 30540 19556 30564 19558
rect 30620 19556 30644 19558
rect 30700 19556 30706 19558
rect 30398 19547 30706 19556
rect 30398 18524 30706 18533
rect 30398 18522 30404 18524
rect 30460 18522 30484 18524
rect 30540 18522 30564 18524
rect 30620 18522 30644 18524
rect 30700 18522 30706 18524
rect 30460 18470 30462 18522
rect 30642 18470 30644 18522
rect 30398 18468 30404 18470
rect 30460 18468 30484 18470
rect 30540 18468 30564 18470
rect 30620 18468 30644 18470
rect 30700 18468 30706 18470
rect 30398 18459 30706 18468
rect 30398 17436 30706 17445
rect 30398 17434 30404 17436
rect 30460 17434 30484 17436
rect 30540 17434 30564 17436
rect 30620 17434 30644 17436
rect 30700 17434 30706 17436
rect 30460 17382 30462 17434
rect 30642 17382 30644 17434
rect 30398 17380 30404 17382
rect 30460 17380 30484 17382
rect 30540 17380 30564 17382
rect 30620 17380 30644 17382
rect 30700 17380 30706 17382
rect 30398 17371 30706 17380
rect 30398 16348 30706 16357
rect 30398 16346 30404 16348
rect 30460 16346 30484 16348
rect 30540 16346 30564 16348
rect 30620 16346 30644 16348
rect 30700 16346 30706 16348
rect 30460 16294 30462 16346
rect 30642 16294 30644 16346
rect 30398 16292 30404 16294
rect 30460 16292 30484 16294
rect 30540 16292 30564 16294
rect 30620 16292 30644 16294
rect 30700 16292 30706 16294
rect 30398 16283 30706 16292
rect 30398 15260 30706 15269
rect 30398 15258 30404 15260
rect 30460 15258 30484 15260
rect 30540 15258 30564 15260
rect 30620 15258 30644 15260
rect 30700 15258 30706 15260
rect 30460 15206 30462 15258
rect 30642 15206 30644 15258
rect 30398 15204 30404 15206
rect 30460 15204 30484 15206
rect 30540 15204 30564 15206
rect 30620 15204 30644 15206
rect 30700 15204 30706 15206
rect 30398 15195 30706 15204
rect 30398 14172 30706 14181
rect 30398 14170 30404 14172
rect 30460 14170 30484 14172
rect 30540 14170 30564 14172
rect 30620 14170 30644 14172
rect 30700 14170 30706 14172
rect 30460 14118 30462 14170
rect 30642 14118 30644 14170
rect 30398 14116 30404 14118
rect 30460 14116 30484 14118
rect 30540 14116 30564 14118
rect 30620 14116 30644 14118
rect 30700 14116 30706 14118
rect 30398 14107 30706 14116
rect 30398 13084 30706 13093
rect 30398 13082 30404 13084
rect 30460 13082 30484 13084
rect 30540 13082 30564 13084
rect 30620 13082 30644 13084
rect 30700 13082 30706 13084
rect 30460 13030 30462 13082
rect 30642 13030 30644 13082
rect 30398 13028 30404 13030
rect 30460 13028 30484 13030
rect 30540 13028 30564 13030
rect 30620 13028 30644 13030
rect 30700 13028 30706 13030
rect 30398 13019 30706 13028
rect 29736 12232 29788 12238
rect 29736 12174 29788 12180
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 29644 3188 29696 3194
rect 29644 3130 29696 3136
rect 28908 3052 28960 3058
rect 28908 2994 28960 3000
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 28816 2440 28868 2446
rect 28920 2428 28948 2994
rect 29748 2514 29776 12174
rect 30840 12096 30892 12102
rect 30840 12038 30892 12044
rect 30398 11996 30706 12005
rect 30398 11994 30404 11996
rect 30460 11994 30484 11996
rect 30540 11994 30564 11996
rect 30620 11994 30644 11996
rect 30700 11994 30706 11996
rect 30460 11942 30462 11994
rect 30642 11942 30644 11994
rect 30398 11940 30404 11942
rect 30460 11940 30484 11942
rect 30540 11940 30564 11942
rect 30620 11940 30644 11942
rect 30700 11940 30706 11942
rect 30398 11931 30706 11940
rect 30852 11898 30880 12038
rect 30840 11892 30892 11898
rect 30840 11834 30892 11840
rect 30398 10908 30706 10917
rect 30398 10906 30404 10908
rect 30460 10906 30484 10908
rect 30540 10906 30564 10908
rect 30620 10906 30644 10908
rect 30700 10906 30706 10908
rect 30460 10854 30462 10906
rect 30642 10854 30644 10906
rect 30398 10852 30404 10854
rect 30460 10852 30484 10854
rect 30540 10852 30564 10854
rect 30620 10852 30644 10854
rect 30700 10852 30706 10854
rect 30398 10843 30706 10852
rect 30944 10742 30972 22066
rect 31128 13190 31156 24686
rect 31312 24274 31340 24686
rect 31300 24268 31352 24274
rect 31300 24210 31352 24216
rect 31312 17746 31340 24210
rect 31404 19334 31432 26710
rect 31482 26616 31538 26625
rect 31482 26551 31484 26560
rect 31536 26551 31538 26560
rect 31484 26522 31536 26528
rect 31772 26518 31800 26846
rect 31760 26512 31812 26518
rect 31760 26454 31812 26460
rect 31852 26512 31904 26518
rect 31852 26454 31904 26460
rect 31576 26444 31628 26450
rect 31576 26386 31628 26392
rect 31668 26444 31720 26450
rect 31668 26386 31720 26392
rect 31588 26353 31616 26386
rect 31574 26344 31630 26353
rect 31574 26279 31630 26288
rect 31680 26042 31708 26386
rect 31864 26353 31892 26454
rect 32048 26353 32076 26930
rect 31850 26344 31906 26353
rect 31760 26308 31812 26314
rect 31850 26279 31906 26288
rect 32034 26344 32090 26353
rect 32034 26279 32090 26288
rect 31760 26250 31812 26256
rect 31772 26042 31800 26250
rect 31668 26036 31720 26042
rect 31668 25978 31720 25984
rect 31760 26036 31812 26042
rect 31760 25978 31812 25984
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31772 24614 31800 24754
rect 31760 24608 31812 24614
rect 31760 24550 31812 24556
rect 31404 19306 31524 19334
rect 31300 17740 31352 17746
rect 31300 17682 31352 17688
rect 31116 13184 31168 13190
rect 31116 13126 31168 13132
rect 30932 10736 30984 10742
rect 30932 10678 30984 10684
rect 30398 9820 30706 9829
rect 30398 9818 30404 9820
rect 30460 9818 30484 9820
rect 30540 9818 30564 9820
rect 30620 9818 30644 9820
rect 30700 9818 30706 9820
rect 30460 9766 30462 9818
rect 30642 9766 30644 9818
rect 30398 9764 30404 9766
rect 30460 9764 30484 9766
rect 30540 9764 30564 9766
rect 30620 9764 30644 9766
rect 30700 9764 30706 9766
rect 30398 9755 30706 9764
rect 30398 8732 30706 8741
rect 30398 8730 30404 8732
rect 30460 8730 30484 8732
rect 30540 8730 30564 8732
rect 30620 8730 30644 8732
rect 30700 8730 30706 8732
rect 30460 8678 30462 8730
rect 30642 8678 30644 8730
rect 30398 8676 30404 8678
rect 30460 8676 30484 8678
rect 30540 8676 30564 8678
rect 30620 8676 30644 8678
rect 30700 8676 30706 8678
rect 30398 8667 30706 8676
rect 30398 7644 30706 7653
rect 30398 7642 30404 7644
rect 30460 7642 30484 7644
rect 30540 7642 30564 7644
rect 30620 7642 30644 7644
rect 30700 7642 30706 7644
rect 30460 7590 30462 7642
rect 30642 7590 30644 7642
rect 30398 7588 30404 7590
rect 30460 7588 30484 7590
rect 30540 7588 30564 7590
rect 30620 7588 30644 7590
rect 30700 7588 30706 7590
rect 30398 7579 30706 7588
rect 30398 6556 30706 6565
rect 30398 6554 30404 6556
rect 30460 6554 30484 6556
rect 30540 6554 30564 6556
rect 30620 6554 30644 6556
rect 30700 6554 30706 6556
rect 30460 6502 30462 6554
rect 30642 6502 30644 6554
rect 30398 6500 30404 6502
rect 30460 6500 30484 6502
rect 30540 6500 30564 6502
rect 30620 6500 30644 6502
rect 30700 6500 30706 6502
rect 30398 6491 30706 6500
rect 30398 5468 30706 5477
rect 30398 5466 30404 5468
rect 30460 5466 30484 5468
rect 30540 5466 30564 5468
rect 30620 5466 30644 5468
rect 30700 5466 30706 5468
rect 30460 5414 30462 5466
rect 30642 5414 30644 5466
rect 30398 5412 30404 5414
rect 30460 5412 30484 5414
rect 30540 5412 30564 5414
rect 30620 5412 30644 5414
rect 30700 5412 30706 5414
rect 30398 5403 30706 5412
rect 30398 4380 30706 4389
rect 30398 4378 30404 4380
rect 30460 4378 30484 4380
rect 30540 4378 30564 4380
rect 30620 4378 30644 4380
rect 30700 4378 30706 4380
rect 30460 4326 30462 4378
rect 30642 4326 30644 4378
rect 30398 4324 30404 4326
rect 30460 4324 30484 4326
rect 30540 4324 30564 4326
rect 30620 4324 30644 4326
rect 30700 4324 30706 4326
rect 30398 4315 30706 4324
rect 31496 3942 31524 19306
rect 31772 9926 31800 24550
rect 32140 12986 32168 26930
rect 32784 15366 32812 27338
rect 32876 27130 32904 29200
rect 33048 27600 33100 27606
rect 33046 27568 33048 27577
rect 33100 27568 33102 27577
rect 33336 27538 33364 29294
rect 33506 29200 33562 29294
rect 34716 29294 34850 29322
rect 34058 27704 34114 27713
rect 34058 27639 34114 27648
rect 33046 27503 33102 27512
rect 33324 27532 33376 27538
rect 33324 27474 33376 27480
rect 33600 27464 33652 27470
rect 33600 27406 33652 27412
rect 33612 27305 33640 27406
rect 33968 27328 34020 27334
rect 33598 27296 33654 27305
rect 33968 27270 34020 27276
rect 33598 27231 33654 27240
rect 32864 27124 32916 27130
rect 32864 27066 32916 27072
rect 33876 27124 33928 27130
rect 33876 27066 33928 27072
rect 33600 26852 33652 26858
rect 33600 26794 33652 26800
rect 33612 26625 33640 26794
rect 33598 26616 33654 26625
rect 33598 26551 33654 26560
rect 33888 26489 33916 27066
rect 33980 27062 34008 27270
rect 33968 27056 34020 27062
rect 33968 26998 34020 27004
rect 34072 26790 34100 27639
rect 34716 27538 34744 29294
rect 34794 29200 34850 29294
rect 35438 29200 35494 30000
rect 36082 29322 36138 30000
rect 36082 29294 36308 29322
rect 36082 29200 36138 29294
rect 34888 27600 34940 27606
rect 34888 27542 34940 27548
rect 34704 27532 34756 27538
rect 34704 27474 34756 27480
rect 34900 27470 34928 27542
rect 34888 27464 34940 27470
rect 34888 27406 34940 27412
rect 35072 27464 35124 27470
rect 35072 27406 35124 27412
rect 35346 27432 35402 27441
rect 34888 27056 34940 27062
rect 34610 27024 34666 27033
rect 34888 26998 34940 27004
rect 34610 26959 34612 26968
rect 34664 26959 34666 26968
rect 34612 26930 34664 26936
rect 34060 26784 34112 26790
rect 34060 26726 34112 26732
rect 33874 26480 33930 26489
rect 33874 26415 33930 26424
rect 34900 26042 34928 26998
rect 34980 26852 35032 26858
rect 34980 26794 35032 26800
rect 34992 26625 35020 26794
rect 34978 26616 35034 26625
rect 34978 26551 35034 26560
rect 34888 26036 34940 26042
rect 34888 25978 34940 25984
rect 32864 25288 32916 25294
rect 32864 25230 32916 25236
rect 32876 24954 32904 25230
rect 34520 25220 34572 25226
rect 34520 25162 34572 25168
rect 32864 24948 32916 24954
rect 32864 24890 32916 24896
rect 32864 24744 32916 24750
rect 32864 24686 32916 24692
rect 32772 15360 32824 15366
rect 32772 15302 32824 15308
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 32324 12442 32352 12786
rect 32312 12436 32364 12442
rect 32876 12434 32904 24686
rect 34532 24410 34560 25162
rect 34520 24404 34572 24410
rect 34520 24346 34572 24352
rect 35084 22094 35112 27406
rect 35346 27367 35402 27376
rect 35254 27024 35310 27033
rect 35254 26959 35310 26968
rect 35162 26616 35218 26625
rect 35162 26551 35218 26560
rect 35176 26246 35204 26551
rect 35164 26240 35216 26246
rect 35164 26182 35216 26188
rect 35268 25906 35296 26959
rect 35360 26246 35388 27367
rect 35452 27130 35480 29200
rect 36280 27402 36308 29294
rect 37370 29200 37426 30000
rect 38014 29322 38070 30000
rect 38014 29294 38148 29322
rect 38014 29200 38070 29294
rect 37384 27470 37412 29200
rect 37372 27464 37424 27470
rect 37372 27406 37424 27412
rect 37922 27432 37978 27441
rect 36268 27396 36320 27402
rect 36268 27338 36320 27344
rect 37648 27396 37700 27402
rect 37922 27367 37924 27376
rect 37648 27338 37700 27344
rect 37976 27367 37978 27376
rect 37924 27338 37976 27344
rect 35808 27328 35860 27334
rect 35860 27288 35940 27316
rect 35808 27270 35860 27276
rect 35440 27124 35492 27130
rect 35440 27066 35492 27072
rect 35716 26988 35768 26994
rect 35452 26948 35716 26976
rect 35348 26240 35400 26246
rect 35348 26182 35400 26188
rect 35256 25900 35308 25906
rect 35256 25842 35308 25848
rect 35452 24138 35480 26948
rect 35716 26930 35768 26936
rect 35808 26988 35860 26994
rect 35808 26930 35860 26936
rect 35820 26489 35848 26930
rect 35806 26480 35862 26489
rect 35912 26450 35940 27288
rect 36636 26988 36688 26994
rect 36636 26930 36688 26936
rect 35806 26415 35808 26424
rect 35860 26415 35862 26424
rect 35900 26444 35952 26450
rect 35808 26386 35860 26392
rect 35900 26386 35952 26392
rect 35532 26376 35584 26382
rect 35584 26324 35756 26330
rect 35532 26318 35756 26324
rect 35544 26314 35756 26318
rect 35544 26308 35768 26314
rect 35544 26302 35716 26308
rect 35716 26250 35768 26256
rect 36648 26042 36676 26930
rect 37660 26246 37688 27338
rect 38120 27130 38148 29294
rect 39302 29200 39358 30000
rect 39946 29200 40002 30000
rect 41234 29322 41290 30000
rect 41234 29294 41368 29322
rect 41234 29200 41290 29294
rect 38290 27840 38346 27849
rect 38290 27775 38346 27784
rect 38200 27600 38252 27606
rect 38200 27542 38252 27548
rect 38212 27130 38240 27542
rect 38304 27402 38332 27775
rect 39212 27464 39264 27470
rect 39316 27452 39344 29200
rect 39580 28008 39632 28014
rect 39580 27950 39632 27956
rect 39672 28008 39724 28014
rect 39672 27950 39724 27956
rect 39264 27424 39344 27452
rect 39212 27406 39264 27412
rect 38292 27396 38344 27402
rect 38292 27338 38344 27344
rect 38476 27328 38528 27334
rect 38476 27270 38528 27276
rect 38568 27328 38620 27334
rect 38568 27270 38620 27276
rect 38108 27124 38160 27130
rect 38108 27066 38160 27072
rect 38200 27124 38252 27130
rect 38200 27066 38252 27072
rect 38384 26988 38436 26994
rect 38384 26930 38436 26936
rect 38396 26625 38424 26930
rect 38382 26616 38438 26625
rect 38382 26551 38438 26560
rect 37648 26240 37700 26246
rect 37648 26182 37700 26188
rect 36636 26036 36688 26042
rect 36636 25978 36688 25984
rect 35440 24132 35492 24138
rect 35440 24074 35492 24080
rect 34992 22066 35112 22094
rect 33324 18760 33376 18766
rect 33324 18702 33376 18708
rect 33336 18290 33364 18702
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 33232 18216 33284 18222
rect 33232 18158 33284 18164
rect 33244 17882 33272 18158
rect 33232 17876 33284 17882
rect 33232 17818 33284 17824
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 32312 12378 32364 12384
rect 32784 12406 32904 12434
rect 31760 9920 31812 9926
rect 31760 9862 31812 9868
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 32128 3528 32180 3534
rect 32128 3470 32180 3476
rect 30398 3292 30706 3301
rect 30398 3290 30404 3292
rect 30460 3290 30484 3292
rect 30540 3290 30564 3292
rect 30620 3290 30644 3292
rect 30700 3290 30706 3292
rect 30460 3238 30462 3290
rect 30642 3238 30644 3290
rect 30398 3236 30404 3238
rect 30460 3236 30484 3238
rect 30540 3236 30564 3238
rect 30620 3236 30644 3238
rect 30700 3236 30706 3238
rect 30398 3227 30706 3236
rect 31576 2848 31628 2854
rect 31576 2790 31628 2796
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 29828 2508 29880 2514
rect 29828 2450 29880 2456
rect 28868 2400 28948 2428
rect 28816 2382 28868 2388
rect 28448 2032 28500 2038
rect 28448 1974 28500 1980
rect 28460 1601 28488 1974
rect 28446 1592 28502 1601
rect 28446 1527 28502 1536
rect 28920 1358 28948 2400
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 28908 1352 28960 1358
rect 28908 1294 28960 1300
rect 29012 800 29040 2382
rect 29656 800 29684 2382
rect 29736 2304 29788 2310
rect 29736 2246 29788 2252
rect 29748 1766 29776 2246
rect 29840 2038 29868 2450
rect 31588 2446 31616 2790
rect 32140 2650 32168 3470
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 32784 2514 32812 12406
rect 32956 10532 33008 10538
rect 32956 10474 33008 10480
rect 32968 3126 32996 10474
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 32956 3120 33008 3126
rect 32956 3062 33008 3068
rect 33612 3058 33640 3538
rect 33796 3534 33824 17478
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 34992 3466 35020 22066
rect 37832 17740 37884 17746
rect 37832 17682 37884 17688
rect 37844 14822 37872 17682
rect 37832 14816 37884 14822
rect 37832 14758 37884 14764
rect 36544 10600 36596 10606
rect 36544 10542 36596 10548
rect 35716 4140 35768 4146
rect 35716 4082 35768 4088
rect 34980 3460 35032 3466
rect 34980 3402 35032 3408
rect 33600 3052 33652 3058
rect 33600 2994 33652 3000
rect 34796 3052 34848 3058
rect 34796 2994 34848 3000
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 32864 2848 32916 2854
rect 32864 2790 32916 2796
rect 32772 2508 32824 2514
rect 32772 2450 32824 2456
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 30748 2304 30800 2310
rect 30748 2246 30800 2252
rect 30398 2204 30706 2213
rect 30398 2202 30404 2204
rect 30460 2202 30484 2204
rect 30540 2202 30564 2204
rect 30620 2202 30644 2204
rect 30700 2202 30706 2204
rect 30460 2150 30462 2202
rect 30642 2150 30644 2202
rect 30398 2148 30404 2150
rect 30460 2148 30484 2150
rect 30540 2148 30564 2150
rect 30620 2148 30644 2150
rect 30700 2148 30706 2150
rect 30398 2139 30706 2148
rect 30760 2038 30788 2246
rect 29828 2032 29880 2038
rect 29828 1974 29880 1980
rect 30748 2032 30800 2038
rect 30748 1974 30800 1980
rect 30746 1864 30802 1873
rect 30746 1799 30802 1808
rect 29736 1760 29788 1766
rect 29736 1702 29788 1708
rect 30760 1494 30788 1799
rect 30748 1488 30800 1494
rect 30748 1430 30800 1436
rect 30944 800 30972 2382
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31668 2304 31720 2310
rect 31668 2246 31720 2252
rect 1398 776 1454 785
rect 1398 711 1454 720
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 31312 762 31340 2246
rect 31680 1986 31708 2246
rect 31404 1958 31708 1986
rect 31404 1902 31432 1958
rect 31392 1896 31444 1902
rect 31392 1838 31444 1844
rect 31576 1896 31628 1902
rect 31576 1838 31628 1844
rect 31588 1737 31616 1838
rect 31574 1728 31630 1737
rect 31574 1663 31630 1672
rect 31668 1488 31720 1494
rect 31668 1430 31720 1436
rect 31680 1290 31708 1430
rect 31668 1284 31720 1290
rect 31668 1226 31720 1232
rect 31496 870 31616 898
rect 31496 762 31524 870
rect 31588 800 31616 870
rect 32876 800 32904 2790
rect 34704 2508 34756 2514
rect 34704 2450 34756 2456
rect 34716 2310 34744 2450
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 34704 2304 34756 2310
rect 34704 2246 34756 2252
rect 33520 800 33548 2246
rect 34808 800 34836 2994
rect 35452 800 35480 2994
rect 35728 2922 35756 4082
rect 36084 3052 36136 3058
rect 36084 2994 36136 3000
rect 35716 2916 35768 2922
rect 35716 2858 35768 2864
rect 36096 800 36124 2994
rect 36268 2848 36320 2854
rect 36268 2790 36320 2796
rect 36280 2446 36308 2790
rect 36268 2440 36320 2446
rect 36268 2382 36320 2388
rect 36556 2378 36584 10542
rect 37648 4480 37700 4486
rect 37648 4422 37700 4428
rect 37660 3058 37688 4422
rect 37648 3052 37700 3058
rect 37648 2994 37700 3000
rect 37844 2990 37872 14758
rect 38488 11898 38516 27270
rect 38580 26489 38608 27270
rect 39592 27146 39620 27950
rect 39684 27334 39712 27950
rect 39960 27606 39988 29200
rect 40868 28076 40920 28082
rect 40868 28018 40920 28024
rect 40408 28008 40460 28014
rect 40222 27976 40278 27985
rect 40408 27950 40460 27956
rect 40222 27911 40278 27920
rect 39948 27600 40000 27606
rect 39948 27542 40000 27548
rect 39672 27328 39724 27334
rect 39672 27270 39724 27276
rect 39856 27328 39908 27334
rect 39856 27270 39908 27276
rect 39592 27118 39712 27146
rect 39684 26926 39712 27118
rect 39868 26994 39896 27270
rect 39856 26988 39908 26994
rect 39856 26930 39908 26936
rect 39304 26920 39356 26926
rect 39304 26862 39356 26868
rect 39672 26920 39724 26926
rect 39672 26862 39724 26868
rect 38566 26480 38622 26489
rect 38566 26415 38622 26424
rect 38476 11892 38528 11898
rect 38476 11834 38528 11840
rect 38476 11552 38528 11558
rect 38476 11494 38528 11500
rect 37740 2984 37792 2990
rect 37740 2926 37792 2932
rect 37832 2984 37884 2990
rect 37832 2926 37884 2932
rect 37648 2848 37700 2854
rect 37648 2790 37700 2796
rect 37660 2446 37688 2790
rect 37648 2440 37700 2446
rect 37648 2382 37700 2388
rect 36544 2372 36596 2378
rect 36544 2314 36596 2320
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 37384 800 37412 2246
rect 37752 2038 37780 2926
rect 37844 2514 37872 2926
rect 38016 2576 38068 2582
rect 38016 2518 38068 2524
rect 37832 2508 37884 2514
rect 37832 2450 37884 2456
rect 37740 2032 37792 2038
rect 37740 1974 37792 1980
rect 38028 800 38056 2518
rect 38488 1902 38516 11494
rect 38568 2576 38620 2582
rect 38568 2518 38620 2524
rect 38476 1896 38528 1902
rect 38580 1873 38608 2518
rect 39316 2446 39344 26862
rect 40236 26246 40264 27911
rect 40420 27538 40448 27950
rect 40880 27946 40908 28018
rect 40868 27940 40920 27946
rect 40868 27882 40920 27888
rect 40960 27940 41012 27946
rect 40960 27882 41012 27888
rect 40592 27600 40644 27606
rect 40684 27600 40736 27606
rect 40592 27542 40644 27548
rect 40682 27568 40684 27577
rect 40736 27568 40738 27577
rect 40408 27532 40460 27538
rect 40408 27474 40460 27480
rect 40604 27470 40632 27542
rect 40682 27503 40738 27512
rect 40500 27464 40552 27470
rect 40500 27406 40552 27412
rect 40592 27464 40644 27470
rect 40592 27406 40644 27412
rect 40314 27160 40370 27169
rect 40512 27130 40540 27406
rect 40868 27328 40920 27334
rect 40868 27270 40920 27276
rect 40314 27095 40316 27104
rect 40368 27095 40370 27104
rect 40500 27124 40552 27130
rect 40316 27066 40368 27072
rect 40500 27066 40552 27072
rect 40776 26444 40828 26450
rect 40776 26386 40828 26392
rect 40224 26240 40276 26246
rect 40224 26182 40276 26188
rect 40788 26081 40816 26386
rect 40774 26072 40830 26081
rect 40774 26007 40830 26016
rect 39396 12368 39448 12374
rect 39396 12310 39448 12316
rect 39408 11694 39436 12310
rect 39396 11688 39448 11694
rect 39396 11630 39448 11636
rect 40132 3664 40184 3670
rect 40132 3606 40184 3612
rect 40314 3632 40370 3641
rect 40038 3088 40094 3097
rect 39580 3052 39632 3058
rect 40038 3023 40094 3032
rect 39580 2994 39632 3000
rect 39396 2848 39448 2854
rect 39396 2790 39448 2796
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 39304 2440 39356 2446
rect 39304 2382 39356 2388
rect 38672 2038 38700 2382
rect 38660 2032 38712 2038
rect 38660 1974 38712 1980
rect 38476 1838 38528 1844
rect 38566 1864 38622 1873
rect 38566 1799 38622 1808
rect 39408 1170 39436 2790
rect 39592 2417 39620 2994
rect 39854 2952 39910 2961
rect 39854 2887 39910 2896
rect 39578 2408 39634 2417
rect 39868 2378 39896 2887
rect 40052 2854 40080 3023
rect 40040 2848 40092 2854
rect 40040 2790 40092 2796
rect 40144 2446 40172 3606
rect 40314 3567 40370 3576
rect 40328 3534 40356 3567
rect 40316 3528 40368 3534
rect 40592 3528 40644 3534
rect 40316 3470 40368 3476
rect 40512 3476 40592 3482
rect 40512 3470 40644 3476
rect 40408 3460 40460 3466
rect 40408 3402 40460 3408
rect 40512 3454 40632 3470
rect 40420 3058 40448 3402
rect 40408 3052 40460 3058
rect 40408 2994 40460 3000
rect 40224 2984 40276 2990
rect 40224 2926 40276 2932
rect 40236 2582 40264 2926
rect 40512 2774 40540 3454
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40512 2746 40632 2774
rect 40224 2576 40276 2582
rect 40224 2518 40276 2524
rect 40132 2440 40184 2446
rect 40132 2382 40184 2388
rect 39578 2343 39634 2352
rect 39856 2372 39908 2378
rect 39856 2314 39908 2320
rect 39948 2304 40000 2310
rect 39948 2246 40000 2252
rect 40500 2304 40552 2310
rect 40500 2246 40552 2252
rect 39316 1142 39436 1170
rect 39316 800 39344 1142
rect 39960 800 39988 2246
rect 40512 1970 40540 2246
rect 40500 1964 40552 1970
rect 40500 1906 40552 1912
rect 40604 800 40632 2746
rect 40696 2582 40724 2926
rect 40684 2576 40736 2582
rect 40684 2518 40736 2524
rect 40880 1970 40908 27270
rect 40972 26761 41000 27882
rect 41236 27532 41288 27538
rect 41236 27474 41288 27480
rect 41248 27010 41276 27474
rect 41340 27130 41368 29294
rect 41878 29200 41934 30000
rect 42522 29322 42578 30000
rect 43810 29322 43866 30000
rect 42522 29294 42748 29322
rect 42522 29200 42578 29294
rect 41420 27940 41472 27946
rect 41420 27882 41472 27888
rect 41432 27402 41460 27882
rect 41892 27470 41920 29200
rect 42720 27588 42748 29294
rect 43810 29294 44128 29322
rect 43810 29200 43866 29294
rect 42800 27600 42852 27606
rect 42720 27560 42800 27588
rect 42800 27542 42852 27548
rect 43810 27568 43866 27577
rect 43810 27503 43812 27512
rect 43864 27503 43866 27512
rect 43812 27474 43864 27480
rect 44100 27470 44128 29294
rect 44454 29200 44510 30000
rect 45742 29322 45798 30000
rect 46386 29322 46442 30000
rect 45742 29294 45876 29322
rect 45742 29200 45798 29294
rect 44468 27470 44496 29200
rect 45122 27772 45430 27781
rect 45122 27770 45128 27772
rect 45184 27770 45208 27772
rect 45264 27770 45288 27772
rect 45344 27770 45368 27772
rect 45424 27770 45430 27772
rect 45184 27718 45186 27770
rect 45366 27718 45368 27770
rect 45122 27716 45128 27718
rect 45184 27716 45208 27718
rect 45264 27716 45288 27718
rect 45344 27716 45368 27718
rect 45424 27716 45430 27718
rect 45122 27707 45430 27716
rect 41880 27464 41932 27470
rect 41880 27406 41932 27412
rect 43352 27464 43404 27470
rect 43352 27406 43404 27412
rect 44088 27464 44140 27470
rect 44088 27406 44140 27412
rect 44456 27464 44508 27470
rect 44456 27406 44508 27412
rect 41420 27396 41472 27402
rect 41420 27338 41472 27344
rect 41512 27328 41564 27334
rect 41972 27328 42024 27334
rect 41564 27288 41644 27316
rect 41512 27270 41564 27276
rect 41616 27130 41644 27288
rect 41972 27270 42024 27276
rect 42616 27328 42668 27334
rect 42616 27270 42668 27276
rect 41878 27160 41934 27169
rect 41328 27124 41380 27130
rect 41328 27066 41380 27072
rect 41604 27124 41656 27130
rect 41878 27095 41934 27104
rect 41604 27066 41656 27072
rect 41892 27062 41920 27095
rect 41880 27056 41932 27062
rect 41248 26982 41368 27010
rect 41236 26920 41288 26926
rect 41236 26862 41288 26868
rect 40958 26752 41014 26761
rect 40958 26687 41014 26696
rect 41142 26616 41198 26625
rect 40960 26580 41012 26586
rect 41248 26586 41276 26862
rect 41142 26551 41198 26560
rect 41236 26580 41288 26586
rect 40960 26522 41012 26528
rect 40972 26489 41000 26522
rect 40958 26480 41014 26489
rect 40958 26415 41014 26424
rect 41052 26376 41104 26382
rect 41156 26364 41184 26551
rect 41236 26522 41288 26528
rect 41236 26444 41288 26450
rect 41236 26386 41288 26392
rect 41104 26336 41184 26364
rect 41248 26353 41276 26386
rect 41234 26344 41290 26353
rect 41052 26318 41104 26324
rect 40960 26308 41012 26314
rect 41234 26279 41290 26288
rect 41340 26330 41368 26982
rect 41420 26988 41472 26994
rect 41616 26982 41828 27010
rect 41880 26998 41932 27004
rect 41616 26976 41644 26982
rect 41472 26948 41644 26976
rect 41420 26930 41472 26936
rect 41696 26920 41748 26926
rect 41696 26862 41748 26868
rect 41340 26314 41460 26330
rect 41340 26308 41472 26314
rect 41340 26302 41420 26308
rect 40960 26250 41012 26256
rect 40972 25906 41000 26250
rect 40960 25900 41012 25906
rect 40960 25842 41012 25848
rect 41340 14958 41368 26302
rect 41420 26250 41472 26256
rect 41708 23202 41736 26862
rect 41800 26353 41828 26982
rect 41786 26344 41842 26353
rect 41786 26279 41842 26288
rect 41524 23174 41736 23202
rect 41328 14952 41380 14958
rect 41328 14894 41380 14900
rect 41340 12374 41368 14894
rect 41328 12368 41380 12374
rect 41328 12310 41380 12316
rect 41524 3534 41552 23174
rect 41984 22094 42012 27270
rect 41708 22066 42012 22094
rect 41512 3528 41564 3534
rect 41512 3470 41564 3476
rect 41234 3224 41290 3233
rect 41234 3159 41236 3168
rect 41288 3159 41290 3168
rect 41236 3130 41288 3136
rect 41708 3058 41736 22066
rect 42524 11552 42576 11558
rect 42524 11494 42576 11500
rect 42536 11218 42564 11494
rect 42524 11212 42576 11218
rect 42524 11154 42576 11160
rect 42628 4622 42656 27270
rect 42708 25288 42760 25294
rect 42708 25230 42760 25236
rect 42720 24682 42748 25230
rect 42708 24676 42760 24682
rect 42708 24618 42760 24624
rect 43364 14890 43392 27406
rect 45848 27130 45876 29294
rect 46386 29294 46704 29322
rect 46386 29200 46442 29294
rect 46480 27940 46532 27946
rect 46480 27882 46532 27888
rect 45926 27160 45982 27169
rect 45652 27124 45704 27130
rect 45652 27066 45704 27072
rect 45836 27124 45888 27130
rect 45926 27095 45982 27104
rect 45836 27066 45888 27072
rect 44088 26852 44140 26858
rect 44088 26794 44140 26800
rect 44100 26625 44128 26794
rect 45122 26684 45430 26693
rect 45122 26682 45128 26684
rect 45184 26682 45208 26684
rect 45264 26682 45288 26684
rect 45344 26682 45368 26684
rect 45424 26682 45430 26684
rect 45184 26630 45186 26682
rect 45366 26630 45368 26682
rect 45122 26628 45128 26630
rect 45184 26628 45208 26630
rect 45264 26628 45288 26630
rect 45344 26628 45368 26630
rect 45424 26628 45430 26630
rect 44086 26616 44142 26625
rect 45122 26619 45430 26628
rect 44086 26551 44142 26560
rect 45664 26518 45692 27066
rect 45940 26858 45968 27095
rect 46492 27062 46520 27882
rect 46572 27396 46624 27402
rect 46572 27338 46624 27344
rect 46584 27062 46612 27338
rect 46480 27056 46532 27062
rect 46480 26998 46532 27004
rect 46572 27056 46624 27062
rect 46572 26998 46624 27004
rect 46204 26988 46256 26994
rect 46204 26930 46256 26936
rect 45928 26852 45980 26858
rect 45928 26794 45980 26800
rect 46216 26586 46244 26930
rect 46584 26586 46612 26998
rect 46204 26580 46256 26586
rect 46204 26522 46256 26528
rect 46572 26580 46624 26586
rect 46572 26522 46624 26528
rect 43444 26512 43496 26518
rect 43442 26480 43444 26489
rect 45652 26512 45704 26518
rect 43496 26480 43498 26489
rect 45652 26454 45704 26460
rect 43442 26415 43498 26424
rect 46676 26382 46704 29294
rect 47030 29200 47086 30000
rect 48318 29200 48374 30000
rect 48962 29322 49018 30000
rect 50250 29322 50306 30000
rect 48962 29294 49280 29322
rect 48962 29200 49018 29294
rect 46756 28076 46808 28082
rect 46756 28018 46808 28024
rect 46768 27402 46796 28018
rect 47044 27418 47072 29200
rect 48332 27470 48360 29200
rect 49148 28008 49200 28014
rect 49148 27950 49200 27956
rect 49054 27840 49110 27849
rect 49054 27775 49110 27784
rect 46756 27396 46808 27402
rect 46756 27338 46808 27344
rect 46860 27390 47072 27418
rect 47216 27464 47268 27470
rect 47216 27406 47268 27412
rect 48320 27464 48372 27470
rect 48320 27406 48372 27412
rect 46860 27334 46888 27390
rect 46848 27328 46900 27334
rect 46848 27270 46900 27276
rect 46848 27056 46900 27062
rect 46848 26998 46900 27004
rect 46756 26580 46808 26586
rect 46756 26522 46808 26528
rect 46664 26376 46716 26382
rect 46664 26318 46716 26324
rect 46768 25906 46796 26522
rect 46860 26314 46888 26998
rect 46940 26784 46992 26790
rect 46940 26726 46992 26732
rect 47124 26784 47176 26790
rect 47124 26726 47176 26732
rect 46848 26308 46900 26314
rect 46848 26250 46900 26256
rect 46756 25900 46808 25906
rect 46756 25842 46808 25848
rect 45122 25596 45430 25605
rect 45122 25594 45128 25596
rect 45184 25594 45208 25596
rect 45264 25594 45288 25596
rect 45344 25594 45368 25596
rect 45424 25594 45430 25596
rect 45184 25542 45186 25594
rect 45366 25542 45368 25594
rect 45122 25540 45128 25542
rect 45184 25540 45208 25542
rect 45264 25540 45288 25542
rect 45344 25540 45368 25542
rect 45424 25540 45430 25542
rect 45122 25531 45430 25540
rect 45122 24508 45430 24517
rect 45122 24506 45128 24508
rect 45184 24506 45208 24508
rect 45264 24506 45288 24508
rect 45344 24506 45368 24508
rect 45424 24506 45430 24508
rect 45184 24454 45186 24506
rect 45366 24454 45368 24506
rect 45122 24452 45128 24454
rect 45184 24452 45208 24454
rect 45264 24452 45288 24454
rect 45344 24452 45368 24454
rect 45424 24452 45430 24454
rect 45122 24443 45430 24452
rect 45122 23420 45430 23429
rect 45122 23418 45128 23420
rect 45184 23418 45208 23420
rect 45264 23418 45288 23420
rect 45344 23418 45368 23420
rect 45424 23418 45430 23420
rect 45184 23366 45186 23418
rect 45366 23366 45368 23418
rect 45122 23364 45128 23366
rect 45184 23364 45208 23366
rect 45264 23364 45288 23366
rect 45344 23364 45368 23366
rect 45424 23364 45430 23366
rect 45122 23355 45430 23364
rect 45122 22332 45430 22341
rect 45122 22330 45128 22332
rect 45184 22330 45208 22332
rect 45264 22330 45288 22332
rect 45344 22330 45368 22332
rect 45424 22330 45430 22332
rect 45184 22278 45186 22330
rect 45366 22278 45368 22330
rect 45122 22276 45128 22278
rect 45184 22276 45208 22278
rect 45264 22276 45288 22278
rect 45344 22276 45368 22278
rect 45424 22276 45430 22278
rect 45122 22267 45430 22276
rect 45122 21244 45430 21253
rect 45122 21242 45128 21244
rect 45184 21242 45208 21244
rect 45264 21242 45288 21244
rect 45344 21242 45368 21244
rect 45424 21242 45430 21244
rect 45184 21190 45186 21242
rect 45366 21190 45368 21242
rect 45122 21188 45128 21190
rect 45184 21188 45208 21190
rect 45264 21188 45288 21190
rect 45344 21188 45368 21190
rect 45424 21188 45430 21190
rect 45122 21179 45430 21188
rect 45122 20156 45430 20165
rect 45122 20154 45128 20156
rect 45184 20154 45208 20156
rect 45264 20154 45288 20156
rect 45344 20154 45368 20156
rect 45424 20154 45430 20156
rect 45184 20102 45186 20154
rect 45366 20102 45368 20154
rect 45122 20100 45128 20102
rect 45184 20100 45208 20102
rect 45264 20100 45288 20102
rect 45344 20100 45368 20102
rect 45424 20100 45430 20102
rect 45122 20091 45430 20100
rect 45122 19068 45430 19077
rect 45122 19066 45128 19068
rect 45184 19066 45208 19068
rect 45264 19066 45288 19068
rect 45344 19066 45368 19068
rect 45424 19066 45430 19068
rect 45184 19014 45186 19066
rect 45366 19014 45368 19066
rect 45122 19012 45128 19014
rect 45184 19012 45208 19014
rect 45264 19012 45288 19014
rect 45344 19012 45368 19014
rect 45424 19012 45430 19014
rect 45122 19003 45430 19012
rect 45122 17980 45430 17989
rect 45122 17978 45128 17980
rect 45184 17978 45208 17980
rect 45264 17978 45288 17980
rect 45344 17978 45368 17980
rect 45424 17978 45430 17980
rect 45184 17926 45186 17978
rect 45366 17926 45368 17978
rect 45122 17924 45128 17926
rect 45184 17924 45208 17926
rect 45264 17924 45288 17926
rect 45344 17924 45368 17926
rect 45424 17924 45430 17926
rect 45122 17915 45430 17924
rect 45122 16892 45430 16901
rect 45122 16890 45128 16892
rect 45184 16890 45208 16892
rect 45264 16890 45288 16892
rect 45344 16890 45368 16892
rect 45424 16890 45430 16892
rect 45184 16838 45186 16890
rect 45366 16838 45368 16890
rect 45122 16836 45128 16838
rect 45184 16836 45208 16838
rect 45264 16836 45288 16838
rect 45344 16836 45368 16838
rect 45424 16836 45430 16838
rect 45122 16827 45430 16836
rect 45122 15804 45430 15813
rect 45122 15802 45128 15804
rect 45184 15802 45208 15804
rect 45264 15802 45288 15804
rect 45344 15802 45368 15804
rect 45424 15802 45430 15804
rect 45184 15750 45186 15802
rect 45366 15750 45368 15802
rect 45122 15748 45128 15750
rect 45184 15748 45208 15750
rect 45264 15748 45288 15750
rect 45344 15748 45368 15750
rect 45424 15748 45430 15750
rect 45122 15739 45430 15748
rect 43352 14884 43404 14890
rect 43352 14826 43404 14832
rect 45122 14716 45430 14725
rect 45122 14714 45128 14716
rect 45184 14714 45208 14716
rect 45264 14714 45288 14716
rect 45344 14714 45368 14716
rect 45424 14714 45430 14716
rect 45184 14662 45186 14714
rect 45366 14662 45368 14714
rect 45122 14660 45128 14662
rect 45184 14660 45208 14662
rect 45264 14660 45288 14662
rect 45344 14660 45368 14662
rect 45424 14660 45430 14662
rect 45122 14651 45430 14660
rect 45122 13628 45430 13637
rect 45122 13626 45128 13628
rect 45184 13626 45208 13628
rect 45264 13626 45288 13628
rect 45344 13626 45368 13628
rect 45424 13626 45430 13628
rect 45184 13574 45186 13626
rect 45366 13574 45368 13626
rect 45122 13572 45128 13574
rect 45184 13572 45208 13574
rect 45264 13572 45288 13574
rect 45344 13572 45368 13574
rect 45424 13572 45430 13574
rect 45122 13563 45430 13572
rect 42984 13252 43036 13258
rect 42984 13194 43036 13200
rect 42616 4616 42668 4622
rect 42616 4558 42668 4564
rect 42432 3528 42484 3534
rect 42430 3496 42432 3505
rect 42484 3496 42486 3505
rect 42430 3431 42486 3440
rect 41788 3392 41840 3398
rect 41788 3334 41840 3340
rect 42432 3392 42484 3398
rect 42432 3334 42484 3340
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 41800 3194 41828 3334
rect 41788 3188 41840 3194
rect 41788 3130 41840 3136
rect 41696 3052 41748 3058
rect 41696 2994 41748 3000
rect 41972 3052 42024 3058
rect 41972 2994 42024 3000
rect 41984 2774 42012 2994
rect 41892 2746 42012 2774
rect 42444 2774 42472 3334
rect 42812 3194 42840 3334
rect 42800 3188 42852 3194
rect 42800 3130 42852 3136
rect 42996 3126 43024 13194
rect 45122 12540 45430 12549
rect 45122 12538 45128 12540
rect 45184 12538 45208 12540
rect 45264 12538 45288 12540
rect 45344 12538 45368 12540
rect 45424 12538 45430 12540
rect 45184 12486 45186 12538
rect 45366 12486 45368 12538
rect 45122 12484 45128 12486
rect 45184 12484 45208 12486
rect 45264 12484 45288 12486
rect 45344 12484 45368 12486
rect 45424 12484 45430 12486
rect 45122 12475 45430 12484
rect 43996 12164 44048 12170
rect 43996 12106 44048 12112
rect 44008 11694 44036 12106
rect 43996 11688 44048 11694
rect 43996 11630 44048 11636
rect 44008 7954 44036 11630
rect 45122 11452 45430 11461
rect 45122 11450 45128 11452
rect 45184 11450 45208 11452
rect 45264 11450 45288 11452
rect 45344 11450 45368 11452
rect 45424 11450 45430 11452
rect 45184 11398 45186 11450
rect 45366 11398 45368 11450
rect 45122 11396 45128 11398
rect 45184 11396 45208 11398
rect 45264 11396 45288 11398
rect 45344 11396 45368 11398
rect 45424 11396 45430 11398
rect 45122 11387 45430 11396
rect 45122 10364 45430 10373
rect 45122 10362 45128 10364
rect 45184 10362 45208 10364
rect 45264 10362 45288 10364
rect 45344 10362 45368 10364
rect 45424 10362 45430 10364
rect 45184 10310 45186 10362
rect 45366 10310 45368 10362
rect 45122 10308 45128 10310
rect 45184 10308 45208 10310
rect 45264 10308 45288 10310
rect 45344 10308 45368 10310
rect 45424 10308 45430 10310
rect 45122 10299 45430 10308
rect 45122 9276 45430 9285
rect 45122 9274 45128 9276
rect 45184 9274 45208 9276
rect 45264 9274 45288 9276
rect 45344 9274 45368 9276
rect 45424 9274 45430 9276
rect 45184 9222 45186 9274
rect 45366 9222 45368 9274
rect 45122 9220 45128 9222
rect 45184 9220 45208 9222
rect 45264 9220 45288 9222
rect 45344 9220 45368 9222
rect 45424 9220 45430 9222
rect 45122 9211 45430 9220
rect 45122 8188 45430 8197
rect 45122 8186 45128 8188
rect 45184 8186 45208 8188
rect 45264 8186 45288 8188
rect 45344 8186 45368 8188
rect 45424 8186 45430 8188
rect 45184 8134 45186 8186
rect 45366 8134 45368 8186
rect 45122 8132 45128 8134
rect 45184 8132 45208 8134
rect 45264 8132 45288 8134
rect 45344 8132 45368 8134
rect 45424 8132 45430 8134
rect 45122 8123 45430 8132
rect 43996 7948 44048 7954
rect 43996 7890 44048 7896
rect 46952 7818 46980 26726
rect 47136 26217 47164 26726
rect 47122 26208 47178 26217
rect 47122 26143 47178 26152
rect 47228 25362 47256 27406
rect 48228 27328 48280 27334
rect 48780 27328 48832 27334
rect 48280 27276 48360 27282
rect 48228 27270 48360 27276
rect 48832 27288 49004 27316
rect 48780 27270 48832 27276
rect 48240 27254 48360 27270
rect 48228 26512 48280 26518
rect 48228 26454 48280 26460
rect 48240 26382 48268 26454
rect 48228 26376 48280 26382
rect 48228 26318 48280 26324
rect 47308 26308 47360 26314
rect 47308 26250 47360 26256
rect 47320 26081 47348 26250
rect 47306 26072 47362 26081
rect 47306 26007 47362 26016
rect 47216 25356 47268 25362
rect 47216 25298 47268 25304
rect 47032 20052 47084 20058
rect 47032 19994 47084 20000
rect 47044 16574 47072 19994
rect 47044 16546 47164 16574
rect 46940 7812 46992 7818
rect 46940 7754 46992 7760
rect 45122 7100 45430 7109
rect 45122 7098 45128 7100
rect 45184 7098 45208 7100
rect 45264 7098 45288 7100
rect 45344 7098 45368 7100
rect 45424 7098 45430 7100
rect 45184 7046 45186 7098
rect 45366 7046 45368 7098
rect 45122 7044 45128 7046
rect 45184 7044 45208 7046
rect 45264 7044 45288 7046
rect 45344 7044 45368 7046
rect 45424 7044 45430 7046
rect 45122 7035 45430 7044
rect 45122 6012 45430 6021
rect 45122 6010 45128 6012
rect 45184 6010 45208 6012
rect 45264 6010 45288 6012
rect 45344 6010 45368 6012
rect 45424 6010 45430 6012
rect 45184 5958 45186 6010
rect 45366 5958 45368 6010
rect 45122 5956 45128 5958
rect 45184 5956 45208 5958
rect 45264 5956 45288 5958
rect 45344 5956 45368 5958
rect 45424 5956 45430 5958
rect 45122 5947 45430 5956
rect 46572 5568 46624 5574
rect 46572 5510 46624 5516
rect 45122 4924 45430 4933
rect 45122 4922 45128 4924
rect 45184 4922 45208 4924
rect 45264 4922 45288 4924
rect 45344 4922 45368 4924
rect 45424 4922 45430 4924
rect 45184 4870 45186 4922
rect 45366 4870 45368 4922
rect 45122 4868 45128 4870
rect 45184 4868 45208 4870
rect 45264 4868 45288 4870
rect 45344 4868 45368 4870
rect 45424 4868 45430 4870
rect 45122 4859 45430 4868
rect 45122 3836 45430 3845
rect 45122 3834 45128 3836
rect 45184 3834 45208 3836
rect 45264 3834 45288 3836
rect 45344 3834 45368 3836
rect 45424 3834 45430 3836
rect 45184 3782 45186 3834
rect 45366 3782 45368 3834
rect 45122 3780 45128 3782
rect 45184 3780 45208 3782
rect 45264 3780 45288 3782
rect 45344 3780 45368 3782
rect 45424 3780 45430 3782
rect 45122 3771 45430 3780
rect 45652 3732 45704 3738
rect 45652 3674 45704 3680
rect 45664 3618 45692 3674
rect 45664 3590 45876 3618
rect 45744 3528 45796 3534
rect 45744 3470 45796 3476
rect 45848 3482 45876 3590
rect 43258 3360 43314 3369
rect 43258 3295 43314 3304
rect 42984 3120 43036 3126
rect 42984 3062 43036 3068
rect 43272 2990 43300 3295
rect 45374 3088 45430 3097
rect 43812 3052 43864 3058
rect 45374 3023 45376 3032
rect 43812 2994 43864 3000
rect 45428 3023 45430 3032
rect 45376 2994 45428 3000
rect 43260 2984 43312 2990
rect 43260 2926 43312 2932
rect 42616 2848 42668 2854
rect 42616 2790 42668 2796
rect 42444 2746 42564 2774
rect 41788 2372 41840 2378
rect 41788 2314 41840 2320
rect 40868 1964 40920 1970
rect 40868 1906 40920 1912
rect 41800 1290 41828 2314
rect 41788 1284 41840 1290
rect 41788 1226 41840 1232
rect 41892 800 41920 2746
rect 42536 800 42564 2746
rect 42628 2514 42656 2790
rect 42616 2508 42668 2514
rect 42616 2450 42668 2456
rect 42708 2440 42760 2446
rect 42708 2382 42760 2388
rect 42720 1834 42748 2382
rect 42708 1828 42760 1834
rect 42708 1770 42760 1776
rect 43824 800 43852 2994
rect 45122 2748 45430 2757
rect 45122 2746 45128 2748
rect 45184 2746 45208 2748
rect 45264 2746 45288 2748
rect 45344 2746 45368 2748
rect 45424 2746 45430 2748
rect 45184 2694 45186 2746
rect 45366 2694 45368 2746
rect 45122 2692 45128 2694
rect 45184 2692 45208 2694
rect 45264 2692 45288 2694
rect 45344 2692 45368 2694
rect 45424 2692 45430 2694
rect 45122 2683 45430 2692
rect 45560 2576 45612 2582
rect 45560 2518 45612 2524
rect 45572 2394 45600 2518
rect 45572 2366 45692 2394
rect 44456 2304 44508 2310
rect 44456 2246 44508 2252
rect 45560 2304 45612 2310
rect 45560 2246 45612 2252
rect 44468 800 44496 2246
rect 45572 1630 45600 2246
rect 45664 1630 45692 2366
rect 45560 1624 45612 1630
rect 45560 1566 45612 1572
rect 45652 1624 45704 1630
rect 45652 1566 45704 1572
rect 45756 800 45784 3470
rect 45848 3454 46336 3482
rect 45836 3392 45888 3398
rect 45836 3334 45888 3340
rect 45848 2990 45876 3334
rect 46202 3224 46258 3233
rect 46202 3159 46258 3168
rect 45836 2984 45888 2990
rect 45836 2926 45888 2932
rect 46216 2854 46244 3159
rect 46308 2854 46336 3454
rect 46388 3052 46440 3058
rect 46388 2994 46440 3000
rect 46204 2848 46256 2854
rect 46204 2790 46256 2796
rect 46296 2848 46348 2854
rect 46296 2790 46348 2796
rect 45928 2440 45980 2446
rect 45928 2382 45980 2388
rect 45940 1834 45968 2382
rect 45928 1828 45980 1834
rect 45928 1770 45980 1776
rect 46400 800 46428 2994
rect 46584 2774 46612 5510
rect 46848 3596 46900 3602
rect 46848 3538 46900 3544
rect 46860 3398 46888 3538
rect 46848 3392 46900 3398
rect 46848 3334 46900 3340
rect 47136 3126 47164 16546
rect 48332 7750 48360 27254
rect 48976 26994 49004 27288
rect 48964 26988 49016 26994
rect 48964 26930 49016 26936
rect 48504 26920 48556 26926
rect 48504 26862 48556 26868
rect 48516 13802 48544 26862
rect 49068 26790 49096 27775
rect 49160 27538 49188 27950
rect 49148 27532 49200 27538
rect 49148 27474 49200 27480
rect 49056 26784 49108 26790
rect 49056 26726 49108 26732
rect 49148 26784 49200 26790
rect 49148 26726 49200 26732
rect 48504 13796 48556 13802
rect 48504 13738 48556 13744
rect 48320 7744 48372 7750
rect 48320 7686 48372 7692
rect 47306 3632 47362 3641
rect 47306 3567 47362 3576
rect 47216 3528 47268 3534
rect 47216 3470 47268 3476
rect 47124 3120 47176 3126
rect 47124 3062 47176 3068
rect 46584 2746 46796 2774
rect 46768 2514 46796 2746
rect 46756 2508 46808 2514
rect 46756 2450 46808 2456
rect 46754 2408 46810 2417
rect 46754 2343 46756 2352
rect 46808 2343 46810 2352
rect 46756 2314 46808 2320
rect 46664 2304 46716 2310
rect 46664 2246 46716 2252
rect 46676 1970 46704 2246
rect 46664 1964 46716 1970
rect 46664 1906 46716 1912
rect 47228 1850 47256 3470
rect 47320 3466 47348 3567
rect 47952 3528 48004 3534
rect 48044 3528 48096 3534
rect 47952 3470 48004 3476
rect 48042 3496 48044 3505
rect 48096 3496 48098 3505
rect 47308 3460 47360 3466
rect 47308 3402 47360 3408
rect 47492 3392 47544 3398
rect 47584 3392 47636 3398
rect 47492 3334 47544 3340
rect 47582 3360 47584 3369
rect 47636 3360 47638 3369
rect 47504 2961 47532 3334
rect 47582 3295 47638 3304
rect 47688 3194 47900 3210
rect 47676 3188 47912 3194
rect 47728 3182 47860 3188
rect 47676 3130 47728 3136
rect 47860 3130 47912 3136
rect 47964 3058 47992 3470
rect 48042 3431 48098 3440
rect 47584 3052 47636 3058
rect 47584 2994 47636 3000
rect 47952 3052 48004 3058
rect 47952 2994 48004 3000
rect 47490 2952 47546 2961
rect 47490 2887 47546 2896
rect 47596 2582 47624 2994
rect 47584 2576 47636 2582
rect 47584 2518 47636 2524
rect 47964 2417 47992 2994
rect 48044 2916 48096 2922
rect 48044 2858 48096 2864
rect 48056 2514 48084 2858
rect 48320 2848 48372 2854
rect 48320 2790 48372 2796
rect 48044 2508 48096 2514
rect 48044 2450 48096 2456
rect 47950 2408 48006 2417
rect 47950 2343 48006 2352
rect 47952 2304 48004 2310
rect 47952 2246 48004 2252
rect 47044 1822 47256 1850
rect 47044 800 47072 1822
rect 47964 1222 47992 2246
rect 47952 1216 48004 1222
rect 47952 1158 48004 1164
rect 48332 800 48360 2790
rect 49160 2446 49188 26726
rect 49252 26382 49280 29294
rect 49988 29294 50306 29322
rect 49700 28008 49752 28014
rect 49700 27950 49752 27956
rect 49240 26376 49292 26382
rect 49240 26318 49292 26324
rect 49712 21690 49740 27950
rect 49988 26858 50016 29294
rect 50250 29200 50306 29294
rect 50894 29322 50950 30000
rect 50894 29294 51028 29322
rect 50894 29200 50950 29294
rect 50804 28144 50856 28150
rect 50804 28086 50856 28092
rect 50712 28076 50764 28082
rect 50712 28018 50764 28024
rect 50252 28008 50304 28014
rect 50252 27950 50304 27956
rect 50264 27577 50292 27950
rect 50528 27600 50580 27606
rect 50250 27568 50306 27577
rect 50250 27503 50306 27512
rect 50434 27568 50490 27577
rect 50528 27542 50580 27548
rect 50434 27503 50490 27512
rect 50160 27464 50212 27470
rect 50160 27406 50212 27412
rect 50068 26988 50120 26994
rect 50068 26930 50120 26936
rect 49976 26852 50028 26858
rect 49976 26794 50028 26800
rect 49976 26240 50028 26246
rect 49976 26182 50028 26188
rect 49988 25906 50016 26182
rect 49976 25900 50028 25906
rect 49976 25842 50028 25848
rect 49700 21684 49752 21690
rect 49700 21626 49752 21632
rect 49884 6792 49936 6798
rect 49884 6734 49936 6740
rect 49896 6458 49924 6734
rect 50080 6662 50108 26930
rect 50172 26858 50200 27406
rect 50252 27328 50304 27334
rect 50448 27305 50476 27503
rect 50252 27270 50304 27276
rect 50434 27296 50490 27305
rect 50160 26852 50212 26858
rect 50160 26794 50212 26800
rect 50172 26489 50200 26794
rect 50158 26480 50214 26489
rect 50158 26415 50214 26424
rect 50158 26344 50214 26353
rect 50158 26279 50214 26288
rect 50172 26246 50200 26279
rect 50160 26240 50212 26246
rect 50264 26228 50292 27270
rect 50434 27231 50490 27240
rect 50344 26988 50396 26994
rect 50344 26930 50396 26936
rect 50356 26382 50384 26930
rect 50540 26625 50568 27542
rect 50620 27396 50672 27402
rect 50620 27338 50672 27344
rect 50632 27305 50660 27338
rect 50618 27296 50674 27305
rect 50618 27231 50674 27240
rect 50724 27062 50752 28018
rect 50816 27878 50844 28086
rect 50804 27872 50856 27878
rect 50804 27814 50856 27820
rect 50896 27872 50948 27878
rect 50896 27814 50948 27820
rect 50908 27169 50936 27814
rect 51000 27334 51028 29294
rect 52182 29200 52238 30000
rect 52826 29322 52882 30000
rect 53470 29322 53526 30000
rect 52826 29294 52960 29322
rect 52826 29200 52882 29294
rect 51814 27568 51870 27577
rect 51814 27503 51870 27512
rect 50988 27328 51040 27334
rect 50988 27270 51040 27276
rect 50894 27160 50950 27169
rect 50894 27095 50950 27104
rect 50620 27056 50672 27062
rect 50620 26998 50672 27004
rect 50712 27056 50764 27062
rect 50712 26998 50764 27004
rect 51172 27056 51224 27062
rect 51172 26998 51224 27004
rect 50632 26761 50660 26998
rect 50712 26920 50764 26926
rect 50712 26862 50764 26868
rect 50618 26752 50674 26761
rect 50618 26687 50674 26696
rect 50526 26616 50582 26625
rect 50526 26551 50582 26560
rect 50724 26489 50752 26862
rect 51184 26840 51212 26998
rect 51724 26920 51776 26926
rect 51724 26862 51776 26868
rect 51092 26812 51212 26840
rect 50896 26580 50948 26586
rect 50896 26522 50948 26528
rect 50804 26512 50856 26518
rect 50710 26480 50766 26489
rect 50804 26454 50856 26460
rect 50710 26415 50766 26424
rect 50344 26376 50396 26382
rect 50344 26318 50396 26324
rect 50528 26240 50580 26246
rect 50264 26200 50528 26228
rect 50160 26182 50212 26188
rect 50528 26182 50580 26188
rect 50816 26042 50844 26454
rect 50908 26217 50936 26522
rect 50986 26344 51042 26353
rect 50986 26279 50988 26288
rect 51040 26279 51042 26288
rect 50988 26250 51040 26256
rect 50894 26208 50950 26217
rect 50894 26143 50950 26152
rect 50804 26036 50856 26042
rect 50804 25978 50856 25984
rect 51092 24290 51120 26812
rect 51632 26784 51684 26790
rect 51170 26752 51226 26761
rect 51632 26726 51684 26732
rect 51170 26687 51226 26696
rect 51184 26586 51212 26687
rect 51262 26616 51318 26625
rect 51172 26580 51224 26586
rect 51262 26551 51318 26560
rect 51172 26522 51224 26528
rect 51276 26314 51304 26551
rect 51448 26512 51500 26518
rect 51448 26454 51500 26460
rect 51264 26308 51316 26314
rect 51264 26250 51316 26256
rect 51092 24262 51212 24290
rect 51080 24200 51132 24206
rect 51080 24142 51132 24148
rect 50712 22092 50764 22098
rect 50712 22034 50764 22040
rect 50620 21888 50672 21894
rect 50620 21830 50672 21836
rect 50528 15020 50580 15026
rect 50528 14962 50580 14968
rect 50436 14476 50488 14482
rect 50436 14418 50488 14424
rect 50068 6656 50120 6662
rect 50068 6598 50120 6604
rect 49884 6452 49936 6458
rect 49884 6394 49936 6400
rect 49700 6316 49752 6322
rect 49700 6258 49752 6264
rect 49148 2440 49200 2446
rect 49148 2382 49200 2388
rect 48964 2304 49016 2310
rect 48964 2246 49016 2252
rect 48976 800 49004 2246
rect 49712 1766 49740 6258
rect 50448 6254 50476 14418
rect 50540 14414 50568 14962
rect 50528 14408 50580 14414
rect 50528 14350 50580 14356
rect 50436 6248 50488 6254
rect 50436 6190 50488 6196
rect 50448 2582 50476 6190
rect 50632 2990 50660 21830
rect 50724 21690 50752 22034
rect 51092 22030 51120 24142
rect 51080 22024 51132 22030
rect 51080 21966 51132 21972
rect 50712 21684 50764 21690
rect 50712 21626 50764 21632
rect 50804 14272 50856 14278
rect 50804 14214 50856 14220
rect 50816 12434 50844 14214
rect 50816 12406 51028 12434
rect 50712 3528 50764 3534
rect 50764 3476 50936 3482
rect 50712 3470 50936 3476
rect 50724 3454 50936 3470
rect 50908 3398 50936 3454
rect 50804 3392 50856 3398
rect 50804 3334 50856 3340
rect 50896 3392 50948 3398
rect 50896 3334 50948 3340
rect 50816 3210 50844 3334
rect 51000 3210 51028 12406
rect 50816 3182 51028 3210
rect 50620 2984 50672 2990
rect 50620 2926 50672 2932
rect 50816 2582 50844 3182
rect 51184 3058 51212 24262
rect 51460 24206 51488 26454
rect 51644 26217 51672 26726
rect 51630 26208 51686 26217
rect 51630 26143 51686 26152
rect 51448 24200 51500 24206
rect 51448 24142 51500 24148
rect 51736 22094 51764 26862
rect 51828 26489 51856 27503
rect 52196 27470 52224 29200
rect 52184 27464 52236 27470
rect 52184 27406 52236 27412
rect 51908 27328 51960 27334
rect 51908 27270 51960 27276
rect 51814 26480 51870 26489
rect 51814 26415 51870 26424
rect 51552 22066 51764 22094
rect 51172 3052 51224 3058
rect 51172 2994 51224 3000
rect 50896 2848 50948 2854
rect 50896 2790 50948 2796
rect 50436 2576 50488 2582
rect 50436 2518 50488 2524
rect 50804 2576 50856 2582
rect 50804 2518 50856 2524
rect 50252 2304 50304 2310
rect 50252 2246 50304 2252
rect 49700 1760 49752 1766
rect 49700 1702 49752 1708
rect 50264 800 50292 2246
rect 50908 800 50936 2790
rect 51552 1834 51580 22066
rect 51632 2372 51684 2378
rect 51632 2314 51684 2320
rect 51540 1828 51592 1834
rect 51540 1770 51592 1776
rect 51644 1766 51672 2314
rect 51920 2310 51948 27270
rect 52932 27130 52960 29294
rect 53470 29294 53788 29322
rect 53470 29200 53526 29294
rect 53104 28144 53156 28150
rect 53104 28086 53156 28092
rect 53010 27296 53066 27305
rect 53010 27231 53066 27240
rect 53024 27130 53052 27231
rect 53116 27169 53144 28086
rect 53472 28008 53524 28014
rect 53472 27950 53524 27956
rect 53484 27606 53512 27950
rect 53472 27600 53524 27606
rect 53286 27568 53342 27577
rect 53472 27542 53524 27548
rect 53286 27503 53342 27512
rect 53196 27328 53248 27334
rect 53194 27296 53196 27305
rect 53248 27296 53250 27305
rect 53194 27231 53250 27240
rect 53102 27160 53158 27169
rect 52920 27124 52972 27130
rect 52920 27066 52972 27072
rect 53012 27124 53064 27130
rect 53102 27095 53158 27104
rect 53012 27066 53064 27072
rect 53300 27062 53328 27503
rect 53288 27056 53340 27062
rect 53288 26998 53340 27004
rect 53760 26382 53788 29294
rect 54758 29200 54814 30000
rect 55402 29200 55458 30000
rect 56690 29200 56746 30000
rect 57334 29200 57390 30000
rect 58622 29322 58678 30000
rect 58622 29294 58756 29322
rect 58622 29200 58678 29294
rect 54668 27872 54720 27878
rect 54668 27814 54720 27820
rect 54116 27600 54168 27606
rect 54116 27542 54168 27548
rect 54024 27396 54076 27402
rect 54024 27338 54076 27344
rect 53840 27328 53892 27334
rect 54036 27305 54064 27338
rect 53840 27270 53892 27276
rect 54022 27296 54078 27305
rect 53852 27062 53880 27270
rect 54022 27231 54078 27240
rect 54024 27124 54076 27130
rect 54024 27066 54076 27072
rect 53840 27056 53892 27062
rect 53840 26998 53892 27004
rect 53932 26920 53984 26926
rect 53932 26862 53984 26868
rect 53748 26376 53800 26382
rect 53392 26314 53604 26330
rect 53748 26318 53800 26324
rect 53380 26308 53616 26314
rect 53432 26302 53564 26308
rect 53380 26250 53432 26256
rect 53564 26250 53616 26256
rect 53840 15564 53892 15570
rect 53840 15506 53892 15512
rect 53852 14822 53880 15506
rect 53840 14816 53892 14822
rect 53840 14758 53892 14764
rect 52184 3528 52236 3534
rect 52184 3470 52236 3476
rect 52000 2508 52052 2514
rect 52000 2450 52052 2456
rect 51816 2304 51868 2310
rect 51816 2246 51868 2252
rect 51908 2304 51960 2310
rect 51908 2246 51960 2252
rect 51828 1766 51856 2246
rect 52012 2145 52040 2450
rect 51998 2136 52054 2145
rect 51998 2071 52054 2080
rect 51632 1760 51684 1766
rect 51632 1702 51684 1708
rect 51816 1760 51868 1766
rect 51816 1702 51868 1708
rect 52012 1630 52040 2071
rect 52000 1624 52052 1630
rect 52000 1566 52052 1572
rect 52196 800 52224 3470
rect 52736 3052 52788 3058
rect 52736 2994 52788 3000
rect 52828 3052 52880 3058
rect 52828 2994 52880 3000
rect 52748 2582 52776 2994
rect 52736 2576 52788 2582
rect 52736 2518 52788 2524
rect 52840 800 52868 2994
rect 52920 2848 52972 2854
rect 52920 2790 52972 2796
rect 52932 2514 52960 2790
rect 52920 2508 52972 2514
rect 52920 2450 52972 2456
rect 53104 2304 53156 2310
rect 53104 2246 53156 2252
rect 53472 2304 53524 2310
rect 53472 2246 53524 2252
rect 53116 1630 53144 2246
rect 53104 1624 53156 1630
rect 53104 1566 53156 1572
rect 53484 800 53512 2246
rect 53852 2145 53880 14758
rect 53944 2446 53972 26862
rect 54036 26858 54064 27066
rect 54024 26852 54076 26858
rect 54024 26794 54076 26800
rect 54128 25906 54156 27542
rect 54680 27538 54708 27814
rect 54484 27532 54536 27538
rect 54668 27532 54720 27538
rect 54536 27492 54616 27520
rect 54484 27474 54536 27480
rect 54300 26920 54352 26926
rect 54300 26862 54352 26868
rect 54312 26790 54340 26862
rect 54300 26784 54352 26790
rect 54300 26726 54352 26732
rect 54392 26784 54444 26790
rect 54392 26726 54444 26732
rect 54404 26450 54432 26726
rect 54392 26444 54444 26450
rect 54392 26386 54444 26392
rect 54484 25968 54536 25974
rect 54484 25910 54536 25916
rect 54116 25900 54168 25906
rect 54116 25842 54168 25848
rect 54496 25430 54524 25910
rect 54484 25424 54536 25430
rect 54484 25366 54536 25372
rect 54484 21548 54536 21554
rect 54484 21490 54536 21496
rect 54496 20942 54524 21490
rect 54588 21010 54616 27492
rect 54668 27474 54720 27480
rect 54772 26518 54800 29200
rect 55312 27328 55364 27334
rect 55310 27296 55312 27305
rect 55364 27296 55366 27305
rect 55310 27231 55366 27240
rect 55128 26988 55180 26994
rect 55128 26930 55180 26936
rect 54760 26512 54812 26518
rect 54760 26454 54812 26460
rect 55140 21078 55168 26930
rect 55128 21072 55180 21078
rect 55128 21014 55180 21020
rect 54576 21004 54628 21010
rect 54576 20946 54628 20952
rect 54484 20936 54536 20942
rect 54484 20878 54536 20884
rect 55324 19334 55352 27231
rect 55416 27130 55444 29200
rect 56704 27452 56732 29200
rect 57058 27840 57114 27849
rect 57058 27775 57114 27784
rect 56520 27424 56732 27452
rect 55680 27328 55732 27334
rect 56416 27328 56468 27334
rect 55680 27270 55732 27276
rect 56414 27296 56416 27305
rect 56468 27296 56470 27305
rect 55404 27124 55456 27130
rect 55404 27066 55456 27072
rect 55692 26994 55720 27270
rect 56414 27231 56470 27240
rect 56520 27130 56548 27424
rect 57072 27402 57100 27775
rect 57348 27418 57376 29200
rect 57612 28076 57664 28082
rect 57612 28018 57664 28024
rect 57060 27396 57112 27402
rect 57348 27390 57560 27418
rect 57060 27338 57112 27344
rect 57532 27130 57560 27390
rect 57624 27334 57652 28018
rect 58360 27526 58572 27554
rect 58360 27470 58388 27526
rect 57704 27464 57756 27470
rect 57704 27406 57756 27412
rect 58164 27464 58216 27470
rect 58164 27406 58216 27412
rect 58348 27464 58400 27470
rect 58348 27406 58400 27412
rect 58440 27464 58492 27470
rect 58440 27406 58492 27412
rect 57612 27328 57664 27334
rect 57716 27305 57744 27406
rect 58072 27396 58124 27402
rect 58072 27338 58124 27344
rect 57612 27270 57664 27276
rect 57702 27296 57758 27305
rect 57702 27231 57758 27240
rect 58084 27130 58112 27338
rect 58176 27282 58204 27406
rect 58176 27254 58296 27282
rect 56508 27124 56560 27130
rect 56508 27066 56560 27072
rect 57520 27124 57572 27130
rect 57520 27066 57572 27072
rect 58072 27124 58124 27130
rect 58072 27066 58124 27072
rect 55496 26988 55548 26994
rect 55680 26988 55732 26994
rect 55548 26948 55628 26976
rect 55496 26930 55548 26936
rect 55600 26874 55628 26948
rect 55680 26930 55732 26936
rect 56324 26988 56376 26994
rect 56324 26930 56376 26936
rect 56692 26988 56744 26994
rect 56692 26930 56744 26936
rect 57336 26988 57388 26994
rect 57336 26930 57388 26936
rect 55864 26920 55916 26926
rect 55600 26868 55864 26874
rect 55600 26862 55916 26868
rect 55600 26846 55904 26862
rect 56336 26518 56364 26930
rect 56324 26512 56376 26518
rect 56324 26454 56376 26460
rect 55680 26240 55732 26246
rect 55680 26182 55732 26188
rect 55692 26042 55720 26182
rect 55680 26036 55732 26042
rect 55680 25978 55732 25984
rect 55496 20936 55548 20942
rect 55496 20878 55548 20884
rect 55324 19306 55444 19334
rect 54576 14952 54628 14958
rect 54576 14894 54628 14900
rect 54588 14414 54616 14894
rect 54576 14408 54628 14414
rect 54576 14350 54628 14356
rect 55416 7562 55444 19306
rect 55508 14618 55536 20878
rect 56704 15502 56732 26930
rect 57244 26920 57296 26926
rect 57244 26862 57296 26868
rect 57256 26761 57284 26862
rect 57242 26752 57298 26761
rect 57242 26687 57298 26696
rect 57348 26518 57376 26930
rect 58268 26926 58296 27254
rect 58072 26920 58124 26926
rect 58072 26862 58124 26868
rect 58256 26920 58308 26926
rect 58256 26862 58308 26868
rect 57336 26512 57388 26518
rect 57336 26454 57388 26460
rect 56876 26376 56928 26382
rect 56876 26318 56928 26324
rect 56784 25832 56836 25838
rect 56784 25774 56836 25780
rect 56692 15496 56744 15502
rect 56692 15438 56744 15444
rect 56140 14952 56192 14958
rect 56140 14894 56192 14900
rect 55496 14612 55548 14618
rect 55496 14554 55548 14560
rect 55508 12238 55536 14554
rect 56152 14074 56180 14894
rect 56140 14068 56192 14074
rect 56140 14010 56192 14016
rect 55496 12232 55548 12238
rect 55496 12174 55548 12180
rect 55416 7534 55536 7562
rect 54116 3120 54168 3126
rect 54116 3062 54168 3068
rect 54024 2576 54076 2582
rect 54024 2518 54076 2524
rect 53932 2440 53984 2446
rect 53932 2382 53984 2388
rect 54036 2378 54064 2518
rect 54128 2446 54156 3062
rect 55404 2848 55456 2854
rect 55404 2790 55456 2796
rect 54116 2440 54168 2446
rect 54116 2382 54168 2388
rect 54760 2440 54812 2446
rect 54760 2382 54812 2388
rect 54024 2372 54076 2378
rect 54024 2314 54076 2320
rect 53838 2136 53894 2145
rect 53838 2071 53894 2080
rect 54772 800 54800 2382
rect 55310 2136 55366 2145
rect 55310 2071 55366 2080
rect 55218 2000 55274 2009
rect 55324 1970 55352 2071
rect 55218 1935 55220 1944
rect 55272 1935 55274 1944
rect 55312 1964 55364 1970
rect 55220 1906 55272 1912
rect 55312 1906 55364 1912
rect 55416 800 55444 2790
rect 55508 2689 55536 7534
rect 56692 3120 56744 3126
rect 56692 3062 56744 3068
rect 55588 3052 55640 3058
rect 55588 2994 55640 3000
rect 55600 2961 55628 2994
rect 55586 2952 55642 2961
rect 55586 2887 55642 2896
rect 56704 2854 56732 3062
rect 55864 2848 55916 2854
rect 55864 2790 55916 2796
rect 56692 2848 56744 2854
rect 56692 2790 56744 2796
rect 55494 2680 55550 2689
rect 55494 2615 55550 2624
rect 55876 2378 55904 2790
rect 56796 2514 56824 25774
rect 56888 25362 56916 26318
rect 58084 25906 58112 26862
rect 58164 26852 58216 26858
rect 58164 26794 58216 26800
rect 58176 25974 58204 26794
rect 58452 26353 58480 27406
rect 58544 27130 58572 27526
rect 58532 27124 58584 27130
rect 58532 27066 58584 27072
rect 58728 26518 58756 29294
rect 59266 29200 59322 30000
rect 59910 29322 59966 30000
rect 59910 29294 60228 29322
rect 59910 29200 59966 29294
rect 59084 28008 59136 28014
rect 59084 27950 59136 27956
rect 59096 27062 59124 27950
rect 59280 27452 59308 29200
rect 59728 27940 59780 27946
rect 59728 27882 59780 27888
rect 59360 27872 59412 27878
rect 59360 27814 59412 27820
rect 59372 27606 59400 27814
rect 59360 27600 59412 27606
rect 59360 27542 59412 27548
rect 59452 27600 59504 27606
rect 59452 27542 59504 27548
rect 59360 27464 59412 27470
rect 59280 27424 59360 27452
rect 59360 27406 59412 27412
rect 59464 27402 59492 27542
rect 59452 27396 59504 27402
rect 59452 27338 59504 27344
rect 59544 27396 59596 27402
rect 59544 27338 59596 27344
rect 59176 27328 59228 27334
rect 59176 27270 59228 27276
rect 59188 27130 59216 27270
rect 59556 27169 59584 27338
rect 59542 27160 59598 27169
rect 59176 27124 59228 27130
rect 59176 27066 59228 27072
rect 59280 27118 59492 27146
rect 59084 27056 59136 27062
rect 59084 26998 59136 27004
rect 59176 26988 59228 26994
rect 59280 26976 59308 27118
rect 59464 27062 59492 27118
rect 59542 27095 59598 27104
rect 59452 27056 59504 27062
rect 59452 26998 59504 27004
rect 59228 26948 59308 26976
rect 59360 26988 59412 26994
rect 59176 26930 59228 26936
rect 59360 26930 59412 26936
rect 59636 26988 59688 26994
rect 59636 26930 59688 26936
rect 59174 26616 59230 26625
rect 59174 26551 59230 26560
rect 58716 26512 58768 26518
rect 58716 26454 58768 26460
rect 58438 26344 58494 26353
rect 59188 26314 59216 26551
rect 58438 26279 58494 26288
rect 59176 26308 59228 26314
rect 59176 26250 59228 26256
rect 58164 25968 58216 25974
rect 58164 25910 58216 25916
rect 58072 25900 58124 25906
rect 58072 25842 58124 25848
rect 58532 25900 58584 25906
rect 58532 25842 58584 25848
rect 58544 25702 58572 25842
rect 57888 25696 57940 25702
rect 57888 25638 57940 25644
rect 58532 25696 58584 25702
rect 58532 25638 58584 25644
rect 56876 25356 56928 25362
rect 56876 25298 56928 25304
rect 57900 25294 57928 25638
rect 57888 25288 57940 25294
rect 57888 25230 57940 25236
rect 58544 14822 58572 25638
rect 59372 19334 59400 26930
rect 59544 26920 59596 26926
rect 59544 26862 59596 26868
rect 59452 25696 59504 25702
rect 59452 25638 59504 25644
rect 59464 25498 59492 25638
rect 59452 25492 59504 25498
rect 59452 25434 59504 25440
rect 59280 19306 59400 19334
rect 58532 14816 58584 14822
rect 58532 14758 58584 14764
rect 57612 13796 57664 13802
rect 57612 13738 57664 13744
rect 57428 5704 57480 5710
rect 57428 5646 57480 5652
rect 57244 4072 57296 4078
rect 57244 4014 57296 4020
rect 57336 4072 57388 4078
rect 57336 4014 57388 4020
rect 56968 3732 57020 3738
rect 56968 3674 57020 3680
rect 57060 3732 57112 3738
rect 57060 3674 57112 3680
rect 56980 3126 57008 3674
rect 57072 3602 57100 3674
rect 57060 3596 57112 3602
rect 57060 3538 57112 3544
rect 57152 3596 57204 3602
rect 57152 3538 57204 3544
rect 57164 3398 57192 3538
rect 57152 3392 57204 3398
rect 57152 3334 57204 3340
rect 57256 3233 57284 4014
rect 57348 3942 57376 4014
rect 57336 3936 57388 3942
rect 57336 3878 57388 3884
rect 57336 3392 57388 3398
rect 57336 3334 57388 3340
rect 57242 3224 57298 3233
rect 57242 3159 57298 3168
rect 56968 3120 57020 3126
rect 56968 3062 57020 3068
rect 57152 3120 57204 3126
rect 57152 3062 57204 3068
rect 56416 2508 56468 2514
rect 56416 2450 56468 2456
rect 56784 2508 56836 2514
rect 56784 2450 56836 2456
rect 55864 2372 55916 2378
rect 55864 2314 55916 2320
rect 55956 2304 56008 2310
rect 55956 2246 56008 2252
rect 55968 1698 55996 2246
rect 56428 1698 56456 2450
rect 56692 2440 56744 2446
rect 56692 2382 56744 2388
rect 55956 1692 56008 1698
rect 55956 1634 56008 1640
rect 56416 1692 56468 1698
rect 56416 1634 56468 1640
rect 56704 800 56732 2382
rect 57164 1154 57192 3062
rect 57152 1148 57204 1154
rect 57152 1090 57204 1096
rect 57348 800 57376 3334
rect 57440 2990 57468 5646
rect 57624 3534 57652 13738
rect 59280 6186 59308 19306
rect 59268 6180 59320 6186
rect 59268 6122 59320 6128
rect 59268 4140 59320 4146
rect 59268 4082 59320 4088
rect 57978 3768 58034 3777
rect 57978 3703 58034 3712
rect 57992 3670 58020 3703
rect 57980 3664 58032 3670
rect 57980 3606 58032 3612
rect 58070 3632 58126 3641
rect 58070 3567 58072 3576
rect 58124 3567 58126 3576
rect 58530 3632 58586 3641
rect 58530 3567 58586 3576
rect 58072 3538 58124 3544
rect 58544 3534 58572 3567
rect 57612 3528 57664 3534
rect 57612 3470 57664 3476
rect 58256 3528 58308 3534
rect 58256 3470 58308 3476
rect 58532 3528 58584 3534
rect 58532 3470 58584 3476
rect 58164 3392 58216 3398
rect 58164 3334 58216 3340
rect 58070 3224 58126 3233
rect 57624 3194 57836 3210
rect 57612 3188 57836 3194
rect 57664 3182 57836 3188
rect 57612 3130 57664 3136
rect 57808 3108 57836 3182
rect 58070 3159 58072 3168
rect 58124 3159 58126 3168
rect 58072 3130 58124 3136
rect 57980 3120 58032 3126
rect 57702 3088 57758 3097
rect 57808 3080 57980 3108
rect 57980 3062 58032 3068
rect 57702 3023 57704 3032
rect 57756 3023 57758 3032
rect 57704 2994 57756 3000
rect 57428 2984 57480 2990
rect 57980 2984 58032 2990
rect 57428 2926 57480 2932
rect 57794 2952 57850 2961
rect 58176 2972 58204 3334
rect 58032 2944 58204 2972
rect 57980 2926 58032 2932
rect 57794 2887 57850 2896
rect 57808 2514 57836 2887
rect 57980 2848 58032 2854
rect 57978 2816 57980 2825
rect 58072 2848 58124 2854
rect 58032 2816 58034 2825
rect 58072 2790 58124 2796
rect 57978 2751 58034 2760
rect 57796 2508 57848 2514
rect 57796 2450 57848 2456
rect 58084 1816 58112 2790
rect 58176 2446 58204 2944
rect 58268 2854 58296 3470
rect 58714 2952 58770 2961
rect 58714 2887 58770 2896
rect 58256 2848 58308 2854
rect 58256 2790 58308 2796
rect 58728 2650 58756 2887
rect 58808 2848 58860 2854
rect 58806 2816 58808 2825
rect 58860 2816 58862 2825
rect 58806 2751 58862 2760
rect 58716 2644 58768 2650
rect 58716 2586 58768 2592
rect 58164 2440 58216 2446
rect 58164 2382 58216 2388
rect 58256 2304 58308 2310
rect 58256 2246 58308 2252
rect 57992 1788 58112 1816
rect 58162 1864 58218 1873
rect 58268 1834 58296 2246
rect 58162 1799 58164 1808
rect 57992 800 58020 1788
rect 58216 1799 58218 1808
rect 58256 1828 58308 1834
rect 58164 1770 58216 1776
rect 58256 1770 58308 1776
rect 58070 1728 58126 1737
rect 58070 1663 58072 1672
rect 58124 1663 58126 1672
rect 58072 1634 58124 1640
rect 59280 800 59308 4082
rect 59360 3936 59412 3942
rect 59360 3878 59412 3884
rect 59372 2378 59400 3878
rect 59556 3466 59584 26862
rect 59648 25945 59676 26930
rect 59740 26625 59768 27882
rect 59846 27228 60154 27237
rect 59846 27226 59852 27228
rect 59908 27226 59932 27228
rect 59988 27226 60012 27228
rect 60068 27226 60092 27228
rect 60148 27226 60154 27228
rect 59908 27174 59910 27226
rect 60090 27174 60092 27226
rect 59846 27172 59852 27174
rect 59908 27172 59932 27174
rect 59988 27172 60012 27174
rect 60068 27172 60092 27174
rect 60148 27172 60154 27174
rect 59846 27163 60154 27172
rect 60200 26994 60228 29294
rect 61198 29200 61254 30000
rect 61842 29200 61898 30000
rect 63130 29322 63186 30000
rect 63774 29322 63830 30000
rect 64418 29322 64474 30000
rect 65706 29322 65762 30000
rect 66350 29322 66406 30000
rect 67638 29322 67694 30000
rect 68282 29322 68338 30000
rect 63130 29294 63264 29322
rect 63130 29200 63186 29294
rect 60646 27704 60702 27713
rect 60646 27639 60702 27648
rect 60830 27704 60886 27713
rect 60830 27639 60886 27648
rect 60280 27464 60332 27470
rect 60280 27406 60332 27412
rect 60188 26988 60240 26994
rect 60188 26930 60240 26936
rect 59726 26616 59782 26625
rect 59726 26551 59782 26560
rect 59846 26140 60154 26149
rect 59846 26138 59852 26140
rect 59908 26138 59932 26140
rect 59988 26138 60012 26140
rect 60068 26138 60092 26140
rect 60148 26138 60154 26140
rect 59908 26086 59910 26138
rect 60090 26086 60092 26138
rect 59846 26084 59852 26086
rect 59908 26084 59932 26086
rect 59988 26084 60012 26086
rect 60068 26084 60092 26086
rect 60148 26084 60154 26086
rect 59846 26075 60154 26084
rect 60292 26042 60320 27406
rect 60660 27402 60688 27639
rect 60740 27532 60792 27538
rect 60740 27474 60792 27480
rect 60648 27396 60700 27402
rect 60648 27338 60700 27344
rect 60752 27169 60780 27474
rect 60844 27334 60872 27639
rect 61212 27606 61240 29200
rect 61476 27940 61528 27946
rect 61476 27882 61528 27888
rect 61108 27600 61160 27606
rect 60922 27568 60978 27577
rect 61108 27542 61160 27548
rect 61200 27600 61252 27606
rect 61200 27542 61252 27548
rect 60922 27503 60924 27512
rect 60976 27503 60978 27512
rect 60924 27474 60976 27480
rect 60832 27328 60884 27334
rect 60832 27270 60884 27276
rect 60922 27296 60978 27305
rect 60922 27231 60978 27240
rect 60738 27160 60794 27169
rect 60738 27095 60794 27104
rect 60384 26982 60596 27010
rect 60384 26761 60412 26982
rect 60464 26920 60516 26926
rect 60464 26862 60516 26868
rect 60370 26752 60426 26761
rect 60370 26687 60426 26696
rect 60476 26246 60504 26862
rect 60568 26858 60596 26982
rect 60556 26852 60608 26858
rect 60556 26794 60608 26800
rect 60648 26784 60700 26790
rect 60554 26752 60610 26761
rect 60936 26772 60964 27231
rect 60648 26726 60700 26732
rect 60752 26744 60964 26772
rect 60554 26687 60610 26696
rect 60568 26586 60596 26687
rect 60556 26580 60608 26586
rect 60556 26522 60608 26528
rect 60554 26480 60610 26489
rect 60554 26415 60610 26424
rect 60568 26246 60596 26415
rect 60660 26353 60688 26726
rect 60646 26344 60702 26353
rect 60752 26314 60780 26744
rect 60922 26616 60978 26625
rect 60922 26551 60978 26560
rect 60646 26279 60702 26288
rect 60740 26308 60792 26314
rect 60740 26250 60792 26256
rect 60464 26240 60516 26246
rect 60464 26182 60516 26188
rect 60556 26240 60608 26246
rect 60556 26182 60608 26188
rect 60280 26036 60332 26042
rect 60280 25978 60332 25984
rect 59634 25936 59690 25945
rect 59634 25871 59690 25880
rect 59648 24614 59676 25871
rect 60372 25832 60424 25838
rect 60372 25774 60424 25780
rect 60384 25702 60412 25774
rect 60936 25770 60964 26551
rect 61120 26382 61148 27542
rect 61200 26852 61252 26858
rect 61200 26794 61252 26800
rect 61212 26489 61240 26794
rect 61488 26790 61516 27882
rect 61750 27568 61806 27577
rect 61750 27503 61806 27512
rect 61764 27470 61792 27503
rect 61752 27464 61804 27470
rect 61752 27406 61804 27412
rect 61856 27418 61884 29200
rect 62948 28008 63000 28014
rect 62948 27950 63000 27956
rect 62120 27872 62172 27878
rect 62120 27814 62172 27820
rect 62132 27538 62160 27814
rect 62120 27532 62172 27538
rect 62120 27474 62172 27480
rect 61856 27390 62160 27418
rect 62132 27334 62160 27390
rect 62120 27328 62172 27334
rect 62120 27270 62172 27276
rect 62302 27160 62358 27169
rect 62358 27118 62620 27146
rect 62302 27095 62358 27104
rect 61752 26988 61804 26994
rect 61752 26930 61804 26936
rect 61936 26988 61988 26994
rect 61936 26930 61988 26936
rect 62316 26982 62528 27010
rect 62592 26994 62620 27118
rect 62960 27062 62988 27950
rect 63236 27538 63264 29294
rect 63774 29294 64184 29322
rect 63774 29200 63830 29294
rect 64156 27538 64184 29294
rect 64418 29294 64828 29322
rect 64418 29200 64474 29294
rect 63224 27532 63276 27538
rect 63224 27474 63276 27480
rect 63316 27532 63368 27538
rect 63316 27474 63368 27480
rect 64144 27532 64196 27538
rect 64144 27474 64196 27480
rect 62948 27056 63000 27062
rect 62948 26998 63000 27004
rect 61476 26784 61528 26790
rect 61476 26726 61528 26732
rect 61764 26586 61792 26930
rect 61948 26790 61976 26930
rect 62212 26920 62264 26926
rect 62316 26908 62344 26982
rect 62264 26880 62344 26908
rect 62396 26920 62448 26926
rect 62212 26862 62264 26868
rect 62396 26862 62448 26868
rect 61844 26784 61896 26790
rect 61844 26726 61896 26732
rect 61936 26784 61988 26790
rect 61936 26726 61988 26732
rect 61752 26580 61804 26586
rect 61752 26522 61804 26528
rect 61198 26480 61254 26489
rect 61198 26415 61254 26424
rect 61750 26480 61806 26489
rect 61750 26415 61752 26424
rect 61804 26415 61806 26424
rect 61752 26386 61804 26392
rect 61016 26376 61068 26382
rect 61016 26318 61068 26324
rect 61108 26376 61160 26382
rect 61108 26318 61160 26324
rect 61028 25770 61056 26318
rect 61856 25906 61884 26726
rect 62224 26353 62252 26862
rect 62302 26752 62358 26761
rect 62408 26738 62436 26862
rect 62500 26761 62528 26982
rect 62580 26988 62632 26994
rect 62580 26930 62632 26936
rect 63224 26784 63276 26790
rect 62358 26710 62436 26738
rect 62486 26752 62542 26761
rect 62302 26687 62358 26696
rect 63224 26726 63276 26732
rect 62486 26687 62542 26696
rect 62210 26344 62266 26353
rect 61936 26308 61988 26314
rect 62210 26279 62266 26288
rect 61936 26250 61988 26256
rect 61844 25900 61896 25906
rect 61844 25842 61896 25848
rect 60924 25764 60976 25770
rect 60924 25706 60976 25712
rect 61016 25764 61068 25770
rect 61016 25706 61068 25712
rect 60372 25696 60424 25702
rect 60372 25638 60424 25644
rect 59846 25052 60154 25061
rect 59846 25050 59852 25052
rect 59908 25050 59932 25052
rect 59988 25050 60012 25052
rect 60068 25050 60092 25052
rect 60148 25050 60154 25052
rect 59908 24998 59910 25050
rect 60090 24998 60092 25050
rect 59846 24996 59852 24998
rect 59908 24996 59932 24998
rect 59988 24996 60012 24998
rect 60068 24996 60092 24998
rect 60148 24996 60154 24998
rect 59846 24987 60154 24996
rect 59636 24608 59688 24614
rect 59636 24550 59688 24556
rect 59846 23964 60154 23973
rect 59846 23962 59852 23964
rect 59908 23962 59932 23964
rect 59988 23962 60012 23964
rect 60068 23962 60092 23964
rect 60148 23962 60154 23964
rect 59908 23910 59910 23962
rect 60090 23910 60092 23962
rect 59846 23908 59852 23910
rect 59908 23908 59932 23910
rect 59988 23908 60012 23910
rect 60068 23908 60092 23910
rect 60148 23908 60154 23910
rect 59846 23899 60154 23908
rect 59846 22876 60154 22885
rect 59846 22874 59852 22876
rect 59908 22874 59932 22876
rect 59988 22874 60012 22876
rect 60068 22874 60092 22876
rect 60148 22874 60154 22876
rect 59908 22822 59910 22874
rect 60090 22822 60092 22874
rect 59846 22820 59852 22822
rect 59908 22820 59932 22822
rect 59988 22820 60012 22822
rect 60068 22820 60092 22822
rect 60148 22820 60154 22822
rect 59846 22811 60154 22820
rect 59846 21788 60154 21797
rect 59846 21786 59852 21788
rect 59908 21786 59932 21788
rect 59988 21786 60012 21788
rect 60068 21786 60092 21788
rect 60148 21786 60154 21788
rect 59908 21734 59910 21786
rect 60090 21734 60092 21786
rect 59846 21732 59852 21734
rect 59908 21732 59932 21734
rect 59988 21732 60012 21734
rect 60068 21732 60092 21734
rect 60148 21732 60154 21734
rect 59846 21723 60154 21732
rect 59846 20700 60154 20709
rect 59846 20698 59852 20700
rect 59908 20698 59932 20700
rect 59988 20698 60012 20700
rect 60068 20698 60092 20700
rect 60148 20698 60154 20700
rect 59908 20646 59910 20698
rect 60090 20646 60092 20698
rect 59846 20644 59852 20646
rect 59908 20644 59932 20646
rect 59988 20644 60012 20646
rect 60068 20644 60092 20646
rect 60148 20644 60154 20646
rect 59846 20635 60154 20644
rect 59846 19612 60154 19621
rect 59846 19610 59852 19612
rect 59908 19610 59932 19612
rect 59988 19610 60012 19612
rect 60068 19610 60092 19612
rect 60148 19610 60154 19612
rect 59908 19558 59910 19610
rect 60090 19558 60092 19610
rect 59846 19556 59852 19558
rect 59908 19556 59932 19558
rect 59988 19556 60012 19558
rect 60068 19556 60092 19558
rect 60148 19556 60154 19558
rect 59846 19547 60154 19556
rect 59846 18524 60154 18533
rect 59846 18522 59852 18524
rect 59908 18522 59932 18524
rect 59988 18522 60012 18524
rect 60068 18522 60092 18524
rect 60148 18522 60154 18524
rect 59908 18470 59910 18522
rect 60090 18470 60092 18522
rect 59846 18468 59852 18470
rect 59908 18468 59932 18470
rect 59988 18468 60012 18470
rect 60068 18468 60092 18470
rect 60148 18468 60154 18470
rect 59846 18459 60154 18468
rect 59846 17436 60154 17445
rect 59846 17434 59852 17436
rect 59908 17434 59932 17436
rect 59988 17434 60012 17436
rect 60068 17434 60092 17436
rect 60148 17434 60154 17436
rect 59908 17382 59910 17434
rect 60090 17382 60092 17434
rect 59846 17380 59852 17382
rect 59908 17380 59932 17382
rect 59988 17380 60012 17382
rect 60068 17380 60092 17382
rect 60148 17380 60154 17382
rect 59846 17371 60154 17380
rect 59728 17332 59780 17338
rect 59728 17274 59780 17280
rect 59636 4140 59688 4146
rect 59636 4082 59688 4088
rect 59648 3942 59676 4082
rect 59636 3936 59688 3942
rect 59636 3878 59688 3884
rect 59634 3768 59690 3777
rect 59634 3703 59636 3712
rect 59688 3703 59690 3712
rect 59636 3674 59688 3680
rect 59544 3460 59596 3466
rect 59544 3402 59596 3408
rect 59556 3126 59584 3402
rect 59544 3120 59596 3126
rect 59544 3062 59596 3068
rect 59740 3058 59768 17274
rect 59846 16348 60154 16357
rect 59846 16346 59852 16348
rect 59908 16346 59932 16348
rect 59988 16346 60012 16348
rect 60068 16346 60092 16348
rect 60148 16346 60154 16348
rect 59908 16294 59910 16346
rect 60090 16294 60092 16346
rect 59846 16292 59852 16294
rect 59908 16292 59932 16294
rect 59988 16292 60012 16294
rect 60068 16292 60092 16294
rect 60148 16292 60154 16294
rect 59846 16283 60154 16292
rect 59846 15260 60154 15269
rect 59846 15258 59852 15260
rect 59908 15258 59932 15260
rect 59988 15258 60012 15260
rect 60068 15258 60092 15260
rect 60148 15258 60154 15260
rect 59908 15206 59910 15258
rect 60090 15206 60092 15258
rect 59846 15204 59852 15206
rect 59908 15204 59932 15206
rect 59988 15204 60012 15206
rect 60068 15204 60092 15206
rect 60148 15204 60154 15206
rect 59846 15195 60154 15204
rect 59846 14172 60154 14181
rect 59846 14170 59852 14172
rect 59908 14170 59932 14172
rect 59988 14170 60012 14172
rect 60068 14170 60092 14172
rect 60148 14170 60154 14172
rect 59908 14118 59910 14170
rect 60090 14118 60092 14170
rect 59846 14116 59852 14118
rect 59908 14116 59932 14118
rect 59988 14116 60012 14118
rect 60068 14116 60092 14118
rect 60148 14116 60154 14118
rect 59846 14107 60154 14116
rect 59846 13084 60154 13093
rect 59846 13082 59852 13084
rect 59908 13082 59932 13084
rect 59988 13082 60012 13084
rect 60068 13082 60092 13084
rect 60148 13082 60154 13084
rect 59908 13030 59910 13082
rect 60090 13030 60092 13082
rect 59846 13028 59852 13030
rect 59908 13028 59932 13030
rect 59988 13028 60012 13030
rect 60068 13028 60092 13030
rect 60148 13028 60154 13030
rect 59846 13019 60154 13028
rect 59846 11996 60154 12005
rect 59846 11994 59852 11996
rect 59908 11994 59932 11996
rect 59988 11994 60012 11996
rect 60068 11994 60092 11996
rect 60148 11994 60154 11996
rect 59908 11942 59910 11994
rect 60090 11942 60092 11994
rect 59846 11940 59852 11942
rect 59908 11940 59932 11942
rect 59988 11940 60012 11942
rect 60068 11940 60092 11942
rect 60148 11940 60154 11942
rect 59846 11931 60154 11940
rect 59846 10908 60154 10917
rect 59846 10906 59852 10908
rect 59908 10906 59932 10908
rect 59988 10906 60012 10908
rect 60068 10906 60092 10908
rect 60148 10906 60154 10908
rect 59908 10854 59910 10906
rect 60090 10854 60092 10906
rect 59846 10852 59852 10854
rect 59908 10852 59932 10854
rect 59988 10852 60012 10854
rect 60068 10852 60092 10854
rect 60148 10852 60154 10854
rect 59846 10843 60154 10852
rect 59846 9820 60154 9829
rect 59846 9818 59852 9820
rect 59908 9818 59932 9820
rect 59988 9818 60012 9820
rect 60068 9818 60092 9820
rect 60148 9818 60154 9820
rect 59908 9766 59910 9818
rect 60090 9766 60092 9818
rect 59846 9764 59852 9766
rect 59908 9764 59932 9766
rect 59988 9764 60012 9766
rect 60068 9764 60092 9766
rect 60148 9764 60154 9766
rect 59846 9755 60154 9764
rect 59846 8732 60154 8741
rect 59846 8730 59852 8732
rect 59908 8730 59932 8732
rect 59988 8730 60012 8732
rect 60068 8730 60092 8732
rect 60148 8730 60154 8732
rect 59908 8678 59910 8730
rect 60090 8678 60092 8730
rect 59846 8676 59852 8678
rect 59908 8676 59932 8678
rect 59988 8676 60012 8678
rect 60068 8676 60092 8678
rect 60148 8676 60154 8678
rect 59846 8667 60154 8676
rect 59846 7644 60154 7653
rect 59846 7642 59852 7644
rect 59908 7642 59932 7644
rect 59988 7642 60012 7644
rect 60068 7642 60092 7644
rect 60148 7642 60154 7644
rect 59908 7590 59910 7642
rect 60090 7590 60092 7642
rect 59846 7588 59852 7590
rect 59908 7588 59932 7590
rect 59988 7588 60012 7590
rect 60068 7588 60092 7590
rect 60148 7588 60154 7590
rect 59846 7579 60154 7588
rect 59846 6556 60154 6565
rect 59846 6554 59852 6556
rect 59908 6554 59932 6556
rect 59988 6554 60012 6556
rect 60068 6554 60092 6556
rect 60148 6554 60154 6556
rect 59908 6502 59910 6554
rect 60090 6502 60092 6554
rect 59846 6500 59852 6502
rect 59908 6500 59932 6502
rect 59988 6500 60012 6502
rect 60068 6500 60092 6502
rect 60148 6500 60154 6502
rect 59846 6491 60154 6500
rect 59846 5468 60154 5477
rect 59846 5466 59852 5468
rect 59908 5466 59932 5468
rect 59988 5466 60012 5468
rect 60068 5466 60092 5468
rect 60148 5466 60154 5468
rect 59908 5414 59910 5466
rect 60090 5414 60092 5466
rect 59846 5412 59852 5414
rect 59908 5412 59932 5414
rect 59988 5412 60012 5414
rect 60068 5412 60092 5414
rect 60148 5412 60154 5414
rect 59846 5403 60154 5412
rect 61016 5024 61068 5030
rect 61016 4966 61068 4972
rect 59846 4380 60154 4389
rect 59846 4378 59852 4380
rect 59908 4378 59932 4380
rect 59988 4378 60012 4380
rect 60068 4378 60092 4380
rect 60148 4378 60154 4380
rect 59908 4326 59910 4378
rect 60090 4326 60092 4378
rect 59846 4324 59852 4326
rect 59908 4324 59932 4326
rect 59988 4324 60012 4326
rect 60068 4324 60092 4326
rect 60148 4324 60154 4326
rect 59846 4315 60154 4324
rect 59820 4140 59872 4146
rect 59820 4082 59872 4088
rect 59832 3670 59860 4082
rect 61028 3670 61056 4966
rect 61752 4208 61804 4214
rect 61752 4150 61804 4156
rect 61764 3942 61792 4150
rect 61752 3936 61804 3942
rect 61752 3878 61804 3884
rect 59820 3664 59872 3670
rect 59820 3606 59872 3612
rect 61016 3664 61068 3670
rect 61016 3606 61068 3612
rect 61660 3596 61712 3602
rect 61660 3538 61712 3544
rect 60280 3460 60332 3466
rect 60280 3402 60332 3408
rect 59846 3292 60154 3301
rect 59846 3290 59852 3292
rect 59908 3290 59932 3292
rect 59988 3290 60012 3292
rect 60068 3290 60092 3292
rect 60148 3290 60154 3292
rect 59908 3238 59910 3290
rect 60090 3238 60092 3290
rect 59846 3236 59852 3238
rect 59908 3236 59932 3238
rect 59988 3236 60012 3238
rect 60068 3236 60092 3238
rect 60148 3236 60154 3238
rect 59846 3227 60154 3236
rect 59728 3052 59780 3058
rect 59728 2994 59780 3000
rect 59452 2984 59504 2990
rect 59452 2926 59504 2932
rect 60004 2984 60056 2990
rect 60004 2926 60056 2932
rect 59464 2650 59492 2926
rect 59452 2644 59504 2650
rect 59452 2586 59504 2592
rect 60016 2582 60044 2926
rect 60004 2576 60056 2582
rect 60004 2518 60056 2524
rect 59360 2372 59412 2378
rect 59360 2314 59412 2320
rect 59846 2204 60154 2213
rect 59846 2202 59852 2204
rect 59908 2202 59932 2204
rect 59988 2202 60012 2204
rect 60068 2202 60092 2204
rect 60148 2202 60154 2204
rect 59908 2150 59910 2202
rect 60090 2150 60092 2202
rect 59846 2148 59852 2150
rect 59908 2148 59932 2150
rect 59988 2148 60012 2150
rect 60068 2148 60092 2150
rect 60148 2148 60154 2150
rect 59846 2139 60154 2148
rect 59924 870 60044 898
rect 59924 800 59952 870
rect 31312 734 31524 762
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60016 762 60044 870
rect 60292 762 60320 3402
rect 61672 3126 61700 3538
rect 61660 3120 61712 3126
rect 61660 3062 61712 3068
rect 61752 3120 61804 3126
rect 61752 3062 61804 3068
rect 61764 2854 61792 3062
rect 61844 3052 61896 3058
rect 61844 2994 61896 3000
rect 61752 2848 61804 2854
rect 60922 2816 60978 2825
rect 61752 2790 61804 2796
rect 60922 2751 60978 2760
rect 60646 2136 60702 2145
rect 60646 2071 60648 2080
rect 60700 2071 60702 2080
rect 60740 2100 60792 2106
rect 60648 2042 60700 2048
rect 60740 2042 60792 2048
rect 60752 1970 60780 2042
rect 60936 2038 60964 2751
rect 61292 2440 61344 2446
rect 61292 2382 61344 2388
rect 61476 2440 61528 2446
rect 61476 2382 61528 2388
rect 61016 2304 61068 2310
rect 61014 2272 61016 2281
rect 61068 2272 61070 2281
rect 61014 2207 61070 2216
rect 60924 2032 60976 2038
rect 61016 2032 61068 2038
rect 60924 1974 60976 1980
rect 61014 2000 61016 2009
rect 61068 2000 61070 2009
rect 60740 1964 60792 1970
rect 60740 1906 60792 1912
rect 60832 1964 60884 1970
rect 61014 1935 61070 1944
rect 60832 1906 60884 1912
rect 60844 1737 60872 1906
rect 61304 1737 61332 2382
rect 60830 1728 60886 1737
rect 60830 1663 60886 1672
rect 61290 1728 61346 1737
rect 61290 1663 61346 1672
rect 61212 870 61332 898
rect 61212 800 61240 870
rect 60016 734 60320 762
rect 61198 0 61254 800
rect 61304 762 61332 870
rect 61488 762 61516 2382
rect 61856 800 61884 2994
rect 61948 2854 61976 26250
rect 63236 26217 63264 26726
rect 63222 26208 63278 26217
rect 63222 26143 63278 26152
rect 63328 26042 63356 27474
rect 63500 27464 63552 27470
rect 64800 27452 64828 29294
rect 65706 29294 66024 29322
rect 65706 29200 65762 29294
rect 64880 27464 64932 27470
rect 64800 27424 64880 27452
rect 63500 27406 63552 27412
rect 64880 27406 64932 27412
rect 65708 27464 65760 27470
rect 65892 27464 65944 27470
rect 65760 27424 65892 27452
rect 65708 27406 65760 27412
rect 65892 27406 65944 27412
rect 63512 26450 63540 27406
rect 64604 27328 64656 27334
rect 64604 27270 64656 27276
rect 64616 26994 64644 27270
rect 65996 26994 66024 29294
rect 66350 29294 66668 29322
rect 66350 29200 66406 29294
rect 66640 27470 66668 29294
rect 67638 29294 68048 29322
rect 67638 29200 67694 29294
rect 68020 27878 68048 29294
rect 68282 29294 68692 29322
rect 68282 29200 68338 29294
rect 68008 27872 68060 27878
rect 68008 27814 68060 27820
rect 66628 27464 66680 27470
rect 66628 27406 66680 27412
rect 66260 27328 66312 27334
rect 66260 27270 66312 27276
rect 68008 27328 68060 27334
rect 68008 27270 68060 27276
rect 68192 27328 68244 27334
rect 68468 27328 68520 27334
rect 68192 27270 68244 27276
rect 68374 27296 68430 27305
rect 63684 26988 63736 26994
rect 64604 26988 64656 26994
rect 63736 26948 64184 26976
rect 63684 26930 63736 26936
rect 64156 26790 64184 26948
rect 64604 26930 64656 26936
rect 64696 26988 64748 26994
rect 64696 26930 64748 26936
rect 65984 26988 66036 26994
rect 65984 26930 66036 26936
rect 64708 26858 64736 26930
rect 64880 26920 64932 26926
rect 64880 26862 64932 26868
rect 64696 26852 64748 26858
rect 64696 26794 64748 26800
rect 64052 26784 64104 26790
rect 64052 26726 64104 26732
rect 64144 26784 64196 26790
rect 64144 26726 64196 26732
rect 63500 26444 63552 26450
rect 63500 26386 63552 26392
rect 63316 26036 63368 26042
rect 63316 25978 63368 25984
rect 64064 25294 64092 26726
rect 64144 25832 64196 25838
rect 64144 25774 64196 25780
rect 64052 25288 64104 25294
rect 64052 25230 64104 25236
rect 64156 15094 64184 25774
rect 64236 25220 64288 25226
rect 64236 25162 64288 25168
rect 64248 24614 64276 25162
rect 64236 24608 64288 24614
rect 64236 24550 64288 24556
rect 64696 15360 64748 15366
rect 64696 15302 64748 15308
rect 64144 15088 64196 15094
rect 64144 15030 64196 15036
rect 64156 14958 64184 15030
rect 64708 15026 64736 15302
rect 64892 15162 64920 26862
rect 66272 26790 66300 27270
rect 66260 26784 66312 26790
rect 66260 26726 66312 26732
rect 65062 26480 65118 26489
rect 65062 26415 65118 26424
rect 64972 15496 65024 15502
rect 64972 15438 65024 15444
rect 64880 15156 64932 15162
rect 64880 15098 64932 15104
rect 64696 15020 64748 15026
rect 64696 14962 64748 14968
rect 64144 14952 64196 14958
rect 64144 14894 64196 14900
rect 63408 11144 63460 11150
rect 63408 11086 63460 11092
rect 61936 2848 61988 2854
rect 61936 2790 61988 2796
rect 62578 2680 62634 2689
rect 62578 2615 62634 2624
rect 62762 2680 62818 2689
rect 62762 2615 62764 2624
rect 62592 2582 62620 2615
rect 62816 2615 62818 2624
rect 62764 2586 62816 2592
rect 62580 2576 62632 2582
rect 62580 2518 62632 2524
rect 63420 2446 63448 11086
rect 64052 3052 64104 3058
rect 64052 2994 64104 3000
rect 64064 2961 64092 2994
rect 64050 2952 64106 2961
rect 64050 2887 64106 2896
rect 63500 2848 63552 2854
rect 63500 2790 63552 2796
rect 63408 2440 63460 2446
rect 63408 2382 63460 2388
rect 63132 2304 63184 2310
rect 63132 2246 63184 2252
rect 63144 800 63172 2246
rect 63512 2038 63540 2790
rect 63776 2644 63828 2650
rect 63776 2586 63828 2592
rect 63500 2032 63552 2038
rect 63500 1974 63552 1980
rect 63788 800 63816 2586
rect 64064 2446 64092 2887
rect 64052 2440 64104 2446
rect 64052 2382 64104 2388
rect 64156 1737 64184 14894
rect 64984 14890 65012 15438
rect 65076 15094 65104 26415
rect 68020 25906 68048 27270
rect 68204 27062 68232 27270
rect 68468 27270 68520 27276
rect 68374 27231 68430 27240
rect 68192 27056 68244 27062
rect 68192 26998 68244 27004
rect 68388 26586 68416 27231
rect 68480 26586 68508 27270
rect 68376 26580 68428 26586
rect 68376 26522 68428 26528
rect 68468 26580 68520 26586
rect 68468 26522 68520 26528
rect 68664 26382 68692 29294
rect 69570 29200 69626 30000
rect 70214 29200 70270 30000
rect 70858 29322 70914 30000
rect 72146 29322 72202 30000
rect 70858 29294 71084 29322
rect 70858 29200 70914 29294
rect 69296 28076 69348 28082
rect 69296 28018 69348 28024
rect 68744 27940 68796 27946
rect 68744 27882 68796 27888
rect 68756 27538 68784 27882
rect 68928 27872 68980 27878
rect 68928 27814 68980 27820
rect 68940 27588 68968 27814
rect 69020 27600 69072 27606
rect 68940 27560 69020 27588
rect 69020 27542 69072 27548
rect 68744 27532 68796 27538
rect 68744 27474 68796 27480
rect 69308 27470 69336 28018
rect 69296 27464 69348 27470
rect 69296 27406 69348 27412
rect 69480 27464 69532 27470
rect 69480 27406 69532 27412
rect 68836 26988 68888 26994
rect 68836 26930 68888 26936
rect 69112 26988 69164 26994
rect 69112 26930 69164 26936
rect 68560 26376 68612 26382
rect 68560 26318 68612 26324
rect 68652 26376 68704 26382
rect 68652 26318 68704 26324
rect 68572 26042 68600 26318
rect 68560 26036 68612 26042
rect 68560 25978 68612 25984
rect 68284 25968 68336 25974
rect 68284 25910 68336 25916
rect 68008 25900 68060 25906
rect 68008 25842 68060 25848
rect 68192 21956 68244 21962
rect 68192 21898 68244 21904
rect 68204 21690 68232 21898
rect 68192 21684 68244 21690
rect 68192 21626 68244 21632
rect 68100 21548 68152 21554
rect 68100 21490 68152 21496
rect 66536 19168 66588 19174
rect 66536 19110 66588 19116
rect 65984 17264 66036 17270
rect 65984 17206 66036 17212
rect 65996 15502 66024 17206
rect 65984 15496 66036 15502
rect 65984 15438 66036 15444
rect 65800 15360 65852 15366
rect 65800 15302 65852 15308
rect 65064 15088 65116 15094
rect 65064 15030 65116 15036
rect 64972 14884 65024 14890
rect 64972 14826 65024 14832
rect 64984 14278 65012 14826
rect 64972 14272 65024 14278
rect 64972 14214 65024 14220
rect 64604 6928 64656 6934
rect 64604 6870 64656 6876
rect 64512 3052 64564 3058
rect 64512 2994 64564 3000
rect 64524 2774 64552 2994
rect 64616 2922 64644 6870
rect 65076 4078 65104 15030
rect 65812 13938 65840 15302
rect 66548 15094 66576 19110
rect 67456 16108 67508 16114
rect 67456 16050 67508 16056
rect 67088 15564 67140 15570
rect 67088 15506 67140 15512
rect 66996 15360 67048 15366
rect 66996 15302 67048 15308
rect 66536 15088 66588 15094
rect 66536 15030 66588 15036
rect 65892 15020 65944 15026
rect 65892 14962 65944 14968
rect 65904 14414 65932 14962
rect 65984 14816 66036 14822
rect 65984 14758 66036 14764
rect 66076 14816 66128 14822
rect 66076 14758 66128 14764
rect 65892 14408 65944 14414
rect 65892 14350 65944 14356
rect 65996 14226 66024 14758
rect 66088 14346 66116 14758
rect 66076 14340 66128 14346
rect 66076 14282 66128 14288
rect 65904 14198 66024 14226
rect 65800 13932 65852 13938
rect 65800 13874 65852 13880
rect 65904 5710 65932 14198
rect 65984 14068 66036 14074
rect 65984 14010 66036 14016
rect 65892 5704 65944 5710
rect 65892 5646 65944 5652
rect 65064 4072 65116 4078
rect 65064 4014 65116 4020
rect 64604 2916 64656 2922
rect 64604 2858 64656 2864
rect 64432 2746 64552 2774
rect 64142 1728 64198 1737
rect 64142 1663 64198 1672
rect 64432 800 64460 2746
rect 65996 2446 66024 14010
rect 66260 13864 66312 13870
rect 66260 13806 66312 13812
rect 66272 12850 66300 13806
rect 67008 12918 67036 15302
rect 67100 14618 67128 15506
rect 67180 15496 67232 15502
rect 67180 15438 67232 15444
rect 67088 14612 67140 14618
rect 67088 14554 67140 14560
rect 66996 12912 67048 12918
rect 66996 12854 67048 12860
rect 66260 12844 66312 12850
rect 66260 12786 66312 12792
rect 66272 10810 66300 12786
rect 67100 12170 67128 14554
rect 67192 14074 67220 15438
rect 67180 14068 67232 14074
rect 67180 14010 67232 14016
rect 67192 12730 67220 14010
rect 67272 12776 67324 12782
rect 67192 12724 67272 12730
rect 67192 12718 67324 12724
rect 67192 12702 67312 12718
rect 67192 12442 67220 12702
rect 67468 12442 67496 16050
rect 67732 15496 67784 15502
rect 67732 15438 67784 15444
rect 67548 15360 67600 15366
rect 67548 15302 67600 15308
rect 67180 12436 67232 12442
rect 67180 12378 67232 12384
rect 67456 12436 67508 12442
rect 67456 12378 67508 12384
rect 67560 12170 67588 15302
rect 67744 13258 67772 15438
rect 67824 14340 67876 14346
rect 67824 14282 67876 14288
rect 67732 13252 67784 13258
rect 67732 13194 67784 13200
rect 67744 12986 67772 13194
rect 67836 12986 67864 14282
rect 67732 12980 67784 12986
rect 67732 12922 67784 12928
rect 67824 12980 67876 12986
rect 67824 12922 67876 12928
rect 67088 12164 67140 12170
rect 67088 12106 67140 12112
rect 67548 12164 67600 12170
rect 67548 12106 67600 12112
rect 66260 10804 66312 10810
rect 66260 10746 66312 10752
rect 66996 3460 67048 3466
rect 66996 3402 67048 3408
rect 66166 3088 66222 3097
rect 67008 3058 67036 3402
rect 66166 3023 66222 3032
rect 66720 3052 66772 3058
rect 66180 2922 66208 3023
rect 66720 2994 66772 3000
rect 66996 3052 67048 3058
rect 66996 2994 67048 3000
rect 66168 2916 66220 2922
rect 66168 2858 66220 2864
rect 66352 2848 66404 2854
rect 66352 2790 66404 2796
rect 65984 2440 66036 2446
rect 65984 2382 66036 2388
rect 66076 2440 66128 2446
rect 66076 2382 66128 2388
rect 65708 2304 65760 2310
rect 65708 2246 65760 2252
rect 65720 800 65748 2246
rect 66088 2106 66116 2382
rect 66076 2100 66128 2106
rect 66076 2042 66128 2048
rect 66364 800 66392 2790
rect 66732 2650 66760 2994
rect 68112 2854 68140 21490
rect 68296 16182 68324 25910
rect 68848 22094 68876 26930
rect 69124 26790 69152 26930
rect 69112 26784 69164 26790
rect 69112 26726 69164 26732
rect 69018 25936 69074 25945
rect 69018 25871 69074 25880
rect 68572 22066 68876 22094
rect 68572 18698 68600 22066
rect 68652 21480 68704 21486
rect 68652 21422 68704 21428
rect 68744 21480 68796 21486
rect 68744 21422 68796 21428
rect 68664 21146 68692 21422
rect 68652 21140 68704 21146
rect 68652 21082 68704 21088
rect 68756 20806 68784 21422
rect 68744 20800 68796 20806
rect 68744 20742 68796 20748
rect 68560 18692 68612 18698
rect 68560 18634 68612 18640
rect 68284 16176 68336 16182
rect 68284 16118 68336 16124
rect 68296 15570 68324 16118
rect 68468 16108 68520 16114
rect 68468 16050 68520 16056
rect 68376 15904 68428 15910
rect 68376 15846 68428 15852
rect 68284 15564 68336 15570
rect 68284 15506 68336 15512
rect 68192 15496 68244 15502
rect 68192 15438 68244 15444
rect 68204 13734 68232 15438
rect 68192 13728 68244 13734
rect 68192 13670 68244 13676
rect 68296 12646 68324 15506
rect 68388 12850 68416 15846
rect 68480 14958 68508 16050
rect 68928 15972 68980 15978
rect 68928 15914 68980 15920
rect 68836 15700 68888 15706
rect 68836 15642 68888 15648
rect 68744 15428 68796 15434
rect 68744 15370 68796 15376
rect 68756 15094 68784 15370
rect 68848 15094 68876 15642
rect 68744 15088 68796 15094
rect 68744 15030 68796 15036
rect 68836 15088 68888 15094
rect 68836 15030 68888 15036
rect 68468 14952 68520 14958
rect 68468 14894 68520 14900
rect 68650 14920 68706 14929
rect 68480 14278 68508 14894
rect 68650 14855 68652 14864
rect 68704 14855 68706 14864
rect 68836 14884 68888 14890
rect 68652 14826 68704 14832
rect 68836 14826 68888 14832
rect 68652 14408 68704 14414
rect 68652 14350 68704 14356
rect 68468 14272 68520 14278
rect 68468 14214 68520 14220
rect 68560 13932 68612 13938
rect 68560 13874 68612 13880
rect 68376 12844 68428 12850
rect 68376 12786 68428 12792
rect 68284 12640 68336 12646
rect 68284 12582 68336 12588
rect 68296 12442 68324 12582
rect 68284 12436 68336 12442
rect 68284 12378 68336 12384
rect 68572 9654 68600 13874
rect 68664 13530 68692 14350
rect 68848 13938 68876 14826
rect 68940 14346 68968 15914
rect 69032 14822 69060 25871
rect 69204 15496 69256 15502
rect 69204 15438 69256 15444
rect 69216 15026 69244 15438
rect 69204 15020 69256 15026
rect 69204 14962 69256 14968
rect 69296 15020 69348 15026
rect 69296 14962 69348 14968
rect 69308 14890 69336 14962
rect 69296 14884 69348 14890
rect 69296 14826 69348 14832
rect 69020 14816 69072 14822
rect 69020 14758 69072 14764
rect 68928 14340 68980 14346
rect 68928 14282 68980 14288
rect 69020 14340 69072 14346
rect 69020 14282 69072 14288
rect 69032 14074 69060 14282
rect 69308 14278 69336 14826
rect 69296 14272 69348 14278
rect 69296 14214 69348 14220
rect 69020 14068 69072 14074
rect 69020 14010 69072 14016
rect 68836 13932 68888 13938
rect 68836 13874 68888 13880
rect 68744 13728 68796 13734
rect 68744 13670 68796 13676
rect 68652 13524 68704 13530
rect 68652 13466 68704 13472
rect 68756 12850 68784 13670
rect 68744 12844 68796 12850
rect 68744 12786 68796 12792
rect 68848 12782 68876 13874
rect 69020 13320 69072 13326
rect 69020 13262 69072 13268
rect 68836 12776 68888 12782
rect 68836 12718 68888 12724
rect 69032 10742 69060 13262
rect 69020 10736 69072 10742
rect 69020 10678 69072 10684
rect 68560 9648 68612 9654
rect 68560 9590 68612 9596
rect 69492 6934 69520 27406
rect 69584 27334 69612 29200
rect 69938 27840 69994 27849
rect 70228 27826 70256 29200
rect 70308 28008 70360 28014
rect 70308 27950 70360 27956
rect 69938 27775 69994 27784
rect 70044 27798 70256 27826
rect 69572 27328 69624 27334
rect 69572 27270 69624 27276
rect 69848 26920 69900 26926
rect 69848 26862 69900 26868
rect 69572 26784 69624 26790
rect 69570 26752 69572 26761
rect 69860 26761 69888 26862
rect 69624 26752 69626 26761
rect 69570 26687 69626 26696
rect 69846 26752 69902 26761
rect 69846 26687 69902 26696
rect 69584 19334 69612 26687
rect 69952 26450 69980 27775
rect 70044 26586 70072 27798
rect 70216 27464 70268 27470
rect 70216 27406 70268 27412
rect 70032 26580 70084 26586
rect 70032 26522 70084 26528
rect 69940 26444 69992 26450
rect 69940 26386 69992 26392
rect 70228 22094 70256 27406
rect 70320 26858 70348 27950
rect 70492 27600 70544 27606
rect 70492 27542 70544 27548
rect 70400 27532 70452 27538
rect 70400 27474 70452 27480
rect 70308 26852 70360 26858
rect 70308 26794 70360 26800
rect 70412 26790 70440 27474
rect 70504 27384 70532 27542
rect 70584 27396 70636 27402
rect 70504 27356 70584 27384
rect 70584 27338 70636 27344
rect 70952 27328 71004 27334
rect 70952 27270 71004 27276
rect 70492 27124 70544 27130
rect 70492 27066 70544 27072
rect 70400 26784 70452 26790
rect 70504 26761 70532 27066
rect 70964 26994 70992 27270
rect 70676 26988 70728 26994
rect 70676 26930 70728 26936
rect 70952 26988 71004 26994
rect 70952 26930 71004 26936
rect 70400 26726 70452 26732
rect 70490 26752 70546 26761
rect 70490 26687 70546 26696
rect 70492 26512 70544 26518
rect 70492 26454 70544 26460
rect 70504 26217 70532 26454
rect 70688 26246 70716 26930
rect 70768 26784 70820 26790
rect 70768 26726 70820 26732
rect 70780 26382 70808 26726
rect 70768 26376 70820 26382
rect 70768 26318 70820 26324
rect 71056 26246 71084 29294
rect 71976 29294 72202 29322
rect 71976 27470 72004 29294
rect 72146 29200 72202 29294
rect 72790 29322 72846 30000
rect 74078 29322 74134 30000
rect 74722 29322 74778 30000
rect 76010 29322 76066 30000
rect 76654 29322 76710 30000
rect 77298 29322 77354 30000
rect 72790 29294 73200 29322
rect 72790 29200 72846 29294
rect 72884 27940 72936 27946
rect 72884 27882 72936 27888
rect 72424 27532 72476 27538
rect 72424 27474 72476 27480
rect 71964 27464 72016 27470
rect 71964 27406 72016 27412
rect 72056 27464 72108 27470
rect 72056 27406 72108 27412
rect 71136 27328 71188 27334
rect 71136 27270 71188 27276
rect 71320 27328 71372 27334
rect 71320 27270 71372 27276
rect 71148 27130 71176 27270
rect 71136 27124 71188 27130
rect 71136 27066 71188 27072
rect 71332 26466 71360 27270
rect 71872 27056 71924 27062
rect 71872 26998 71924 27004
rect 71884 26858 71912 26998
rect 71872 26852 71924 26858
rect 71872 26794 71924 26800
rect 71240 26438 71360 26466
rect 70676 26240 70728 26246
rect 70490 26208 70546 26217
rect 70676 26182 70728 26188
rect 71044 26240 71096 26246
rect 71044 26182 71096 26188
rect 70490 26143 70546 26152
rect 71240 22982 71268 26438
rect 71780 26376 71832 26382
rect 71780 26318 71832 26324
rect 71320 26308 71372 26314
rect 71320 26250 71372 26256
rect 71596 26308 71648 26314
rect 71596 26250 71648 26256
rect 71332 25974 71360 26250
rect 71320 25968 71372 25974
rect 71320 25910 71372 25916
rect 71228 22976 71280 22982
rect 71228 22918 71280 22924
rect 70136 22066 70256 22094
rect 69584 19306 69704 19334
rect 69572 16108 69624 16114
rect 69572 16050 69624 16056
rect 69584 15706 69612 16050
rect 69572 15700 69624 15706
rect 69572 15642 69624 15648
rect 69676 15586 69704 19306
rect 70136 17338 70164 22066
rect 70124 17332 70176 17338
rect 70124 17274 70176 17280
rect 70584 16584 70636 16590
rect 70584 16526 70636 16532
rect 70596 15910 70624 16526
rect 70768 16516 70820 16522
rect 70768 16458 70820 16464
rect 70584 15904 70636 15910
rect 70584 15846 70636 15852
rect 69584 15558 69704 15586
rect 69584 13870 69612 15558
rect 69664 15428 69716 15434
rect 69664 15370 69716 15376
rect 69676 15094 69704 15370
rect 69756 15360 69808 15366
rect 69756 15302 69808 15308
rect 69664 15088 69716 15094
rect 69664 15030 69716 15036
rect 69664 14476 69716 14482
rect 69664 14418 69716 14424
rect 69676 14006 69704 14418
rect 69768 14006 69796 15302
rect 70596 15094 70624 15846
rect 70780 15706 70808 16458
rect 70768 15700 70820 15706
rect 70768 15642 70820 15648
rect 71320 15564 71372 15570
rect 71320 15506 71372 15512
rect 71136 15360 71188 15366
rect 71136 15302 71188 15308
rect 70584 15088 70636 15094
rect 70584 15030 70636 15036
rect 70400 15020 70452 15026
rect 70400 14962 70452 14968
rect 70032 14952 70084 14958
rect 70032 14894 70084 14900
rect 70214 14920 70270 14929
rect 69848 14816 69900 14822
rect 69900 14776 69980 14804
rect 69848 14758 69900 14764
rect 69848 14544 69900 14550
rect 69848 14486 69900 14492
rect 69664 14000 69716 14006
rect 69664 13942 69716 13948
rect 69756 14000 69808 14006
rect 69756 13942 69808 13948
rect 69860 13870 69888 14486
rect 69572 13864 69624 13870
rect 69572 13806 69624 13812
rect 69848 13864 69900 13870
rect 69848 13806 69900 13812
rect 69848 13728 69900 13734
rect 69848 13670 69900 13676
rect 69860 13326 69888 13670
rect 69848 13320 69900 13326
rect 69848 13262 69900 13268
rect 69480 6928 69532 6934
rect 69480 6870 69532 6876
rect 68468 3528 68520 3534
rect 68468 3470 68520 3476
rect 68284 3052 68336 3058
rect 68284 2994 68336 3000
rect 68100 2848 68152 2854
rect 68100 2790 68152 2796
rect 67270 2680 67326 2689
rect 66720 2644 66772 2650
rect 67270 2615 67326 2624
rect 66720 2586 66772 2592
rect 67284 2378 67312 2615
rect 67456 2576 67508 2582
rect 67456 2518 67508 2524
rect 67364 2440 67416 2446
rect 67364 2382 67416 2388
rect 66812 2372 66864 2378
rect 66812 2314 66864 2320
rect 67272 2372 67324 2378
rect 67272 2314 67324 2320
rect 66824 2106 66852 2314
rect 67180 2304 67232 2310
rect 67180 2246 67232 2252
rect 67192 2106 67220 2246
rect 66812 2100 66864 2106
rect 66812 2042 66864 2048
rect 67180 2100 67232 2106
rect 67180 2042 67232 2048
rect 67376 1873 67404 2382
rect 67468 2145 67496 2518
rect 67640 2304 67692 2310
rect 67640 2246 67692 2252
rect 67454 2136 67510 2145
rect 67454 2071 67510 2080
rect 67362 1864 67418 1873
rect 67362 1799 67418 1808
rect 66902 1728 66958 1737
rect 66902 1663 66904 1672
rect 66956 1663 66958 1672
rect 66904 1634 66956 1640
rect 67652 800 67680 2246
rect 68296 800 68324 2994
rect 68480 2922 68508 3470
rect 69572 3052 69624 3058
rect 69572 2994 69624 3000
rect 68468 2916 68520 2922
rect 68468 2858 68520 2864
rect 68928 2576 68980 2582
rect 68928 2518 68980 2524
rect 68940 2310 68968 2518
rect 68928 2304 68980 2310
rect 68928 2246 68980 2252
rect 69584 800 69612 2994
rect 69952 2990 69980 14776
rect 70044 13530 70072 14894
rect 70214 14855 70216 14864
rect 70268 14855 70270 14864
rect 70216 14826 70268 14832
rect 70308 14816 70360 14822
rect 70308 14758 70360 14764
rect 70032 13524 70084 13530
rect 70032 13466 70084 13472
rect 70320 12918 70348 14758
rect 70412 14278 70440 14962
rect 70584 14816 70636 14822
rect 70584 14758 70636 14764
rect 70596 14346 70624 14758
rect 71044 14408 71096 14414
rect 71044 14350 71096 14356
rect 70584 14340 70636 14346
rect 70584 14282 70636 14288
rect 70676 14340 70728 14346
rect 70676 14282 70728 14288
rect 70400 14272 70452 14278
rect 70400 14214 70452 14220
rect 70412 13802 70440 14214
rect 70688 13938 70716 14282
rect 70676 13932 70728 13938
rect 70676 13874 70728 13880
rect 70400 13796 70452 13802
rect 70400 13738 70452 13744
rect 70308 12912 70360 12918
rect 70308 12854 70360 12860
rect 70492 7540 70544 7546
rect 70492 7482 70544 7488
rect 70216 3392 70268 3398
rect 70216 3334 70268 3340
rect 69940 2984 69992 2990
rect 69940 2926 69992 2932
rect 69664 2848 69716 2854
rect 69664 2790 69716 2796
rect 69676 2446 69704 2790
rect 69940 2508 69992 2514
rect 69940 2450 69992 2456
rect 69664 2440 69716 2446
rect 69664 2382 69716 2388
rect 69952 2281 69980 2450
rect 69938 2272 69994 2281
rect 69938 2207 69994 2216
rect 70228 800 70256 3334
rect 70308 3120 70360 3126
rect 70306 3088 70308 3097
rect 70360 3088 70362 3097
rect 70306 3023 70362 3032
rect 70400 3052 70452 3058
rect 70400 2994 70452 3000
rect 70412 2582 70440 2994
rect 70504 2774 70532 7482
rect 70584 4480 70636 4486
rect 70584 4422 70636 4428
rect 70596 3126 70624 4422
rect 70584 3120 70636 3126
rect 70584 3062 70636 3068
rect 70504 2746 70624 2774
rect 70400 2576 70452 2582
rect 70400 2518 70452 2524
rect 70596 2446 70624 2746
rect 70584 2440 70636 2446
rect 70584 2382 70636 2388
rect 70688 2281 70716 13874
rect 70768 13864 70820 13870
rect 70768 13806 70820 13812
rect 70780 12238 70808 13806
rect 71056 12986 71084 14350
rect 71044 12980 71096 12986
rect 71044 12922 71096 12928
rect 70768 12232 70820 12238
rect 70768 12174 70820 12180
rect 70768 3528 70820 3534
rect 70768 3470 70820 3476
rect 70780 2650 70808 3470
rect 70860 3392 70912 3398
rect 70860 3334 70912 3340
rect 70768 2644 70820 2650
rect 70768 2586 70820 2592
rect 70674 2272 70730 2281
rect 70674 2207 70730 2216
rect 70872 800 70900 3334
rect 71148 2378 71176 15302
rect 71228 15088 71280 15094
rect 71228 15030 71280 15036
rect 71240 2922 71268 15030
rect 71332 7546 71360 15506
rect 71412 14544 71464 14550
rect 71412 14486 71464 14492
rect 71424 14074 71452 14486
rect 71504 14408 71556 14414
rect 71504 14350 71556 14356
rect 71412 14068 71464 14074
rect 71412 14010 71464 14016
rect 71516 13938 71544 14350
rect 71504 13932 71556 13938
rect 71504 13874 71556 13880
rect 71412 12096 71464 12102
rect 71412 12038 71464 12044
rect 71320 7540 71372 7546
rect 71320 7482 71372 7488
rect 71424 4486 71452 12038
rect 71412 4480 71464 4486
rect 71412 4422 71464 4428
rect 71608 3534 71636 26250
rect 71792 26246 71820 26318
rect 71780 26240 71832 26246
rect 71872 26240 71924 26246
rect 71780 26182 71832 26188
rect 71870 26208 71872 26217
rect 71924 26208 71926 26217
rect 71870 26143 71926 26152
rect 72068 26042 72096 27406
rect 72436 27305 72464 27474
rect 72422 27296 72478 27305
rect 72422 27231 72478 27240
rect 72608 26988 72660 26994
rect 72608 26930 72660 26936
rect 72516 26784 72568 26790
rect 72516 26726 72568 26732
rect 72238 26616 72294 26625
rect 72238 26551 72294 26560
rect 72252 26450 72280 26551
rect 72240 26444 72292 26450
rect 72240 26386 72292 26392
rect 72056 26036 72108 26042
rect 72056 25978 72108 25984
rect 72528 25945 72556 26726
rect 72514 25936 72570 25945
rect 72514 25871 72570 25880
rect 71872 20800 71924 20806
rect 71872 20742 71924 20748
rect 71884 20466 71912 20742
rect 71872 20460 71924 20466
rect 71872 20402 71924 20408
rect 72056 20256 72108 20262
rect 72056 20198 72108 20204
rect 72068 19854 72096 20198
rect 72056 19848 72108 19854
rect 72056 19790 72108 19796
rect 71688 12232 71740 12238
rect 71688 12174 71740 12180
rect 71700 11762 71728 12174
rect 71688 11756 71740 11762
rect 71688 11698 71740 11704
rect 72620 4078 72648 26930
rect 72700 26784 72752 26790
rect 72700 26726 72752 26732
rect 72712 20942 72740 26726
rect 72792 26308 72844 26314
rect 72792 26250 72844 26256
rect 72804 25906 72832 26250
rect 72792 25900 72844 25906
rect 72792 25842 72844 25848
rect 72896 21010 72924 27882
rect 73172 26994 73200 29294
rect 74078 29294 74488 29322
rect 74078 29200 74134 29294
rect 74460 27878 74488 29294
rect 74722 29294 75132 29322
rect 74722 29200 74778 29294
rect 75000 28008 75052 28014
rect 74906 27976 74962 27985
rect 75000 27950 75052 27956
rect 74906 27911 74962 27920
rect 74448 27872 74500 27878
rect 73802 27840 73858 27849
rect 74448 27814 74500 27820
rect 73802 27775 73858 27784
rect 73160 26988 73212 26994
rect 73160 26930 73212 26936
rect 73068 26784 73120 26790
rect 73066 26752 73068 26761
rect 73120 26752 73122 26761
rect 73066 26687 73122 26696
rect 72884 21004 72936 21010
rect 72884 20946 72936 20952
rect 72700 20936 72752 20942
rect 72700 20878 72752 20884
rect 72792 20800 72844 20806
rect 72792 20742 72844 20748
rect 72804 16574 72832 20742
rect 72804 16546 72924 16574
rect 72608 4072 72660 4078
rect 72608 4014 72660 4020
rect 72332 3732 72384 3738
rect 72332 3674 72384 3680
rect 72240 3664 72292 3670
rect 72240 3606 72292 3612
rect 71596 3528 71648 3534
rect 71596 3470 71648 3476
rect 72148 3528 72200 3534
rect 72148 3470 72200 3476
rect 72056 3392 72108 3398
rect 72056 3334 72108 3340
rect 71320 3052 71372 3058
rect 71320 2994 71372 3000
rect 71228 2916 71280 2922
rect 71228 2858 71280 2864
rect 71240 2446 71268 2858
rect 71332 2650 71360 2994
rect 71320 2644 71372 2650
rect 71320 2586 71372 2592
rect 72068 2514 72096 3334
rect 71872 2508 71924 2514
rect 71872 2450 71924 2456
rect 72056 2508 72108 2514
rect 72056 2450 72108 2456
rect 71228 2440 71280 2446
rect 71228 2382 71280 2388
rect 71320 2440 71372 2446
rect 71320 2382 71372 2388
rect 71044 2372 71096 2378
rect 71044 2314 71096 2320
rect 71136 2372 71188 2378
rect 71136 2314 71188 2320
rect 71056 1902 71084 2314
rect 70952 1896 71004 1902
rect 70950 1864 70952 1873
rect 71044 1896 71096 1902
rect 71004 1864 71006 1873
rect 71044 1838 71096 1844
rect 70950 1799 71006 1808
rect 71332 1698 71360 2382
rect 71884 1698 71912 2450
rect 71320 1692 71372 1698
rect 71320 1634 71372 1640
rect 71872 1692 71924 1698
rect 71872 1634 71924 1640
rect 72160 800 72188 3470
rect 72252 3058 72280 3606
rect 72344 3058 72372 3674
rect 72240 3052 72292 3058
rect 72240 2994 72292 3000
rect 72332 3052 72384 3058
rect 72332 2994 72384 3000
rect 72332 2916 72384 2922
rect 72332 2858 72384 2864
rect 72344 2650 72372 2858
rect 72332 2644 72384 2650
rect 72332 2586 72384 2592
rect 72344 2009 72372 2586
rect 72330 2000 72386 2009
rect 72330 1935 72386 1944
rect 72896 1737 72924 16546
rect 73816 12986 73844 27775
rect 74570 27772 74878 27781
rect 74570 27770 74576 27772
rect 74632 27770 74656 27772
rect 74712 27770 74736 27772
rect 74792 27770 74816 27772
rect 74872 27770 74878 27772
rect 74632 27718 74634 27770
rect 74814 27718 74816 27770
rect 74570 27716 74576 27718
rect 74632 27716 74656 27718
rect 74712 27716 74736 27718
rect 74792 27716 74816 27718
rect 74872 27716 74878 27718
rect 74262 27704 74318 27713
rect 74570 27707 74878 27716
rect 74262 27639 74318 27648
rect 74276 27334 74304 27639
rect 74632 27600 74684 27606
rect 74460 27560 74632 27588
rect 74264 27328 74316 27334
rect 74264 27270 74316 27276
rect 74460 26994 74488 27560
rect 74632 27542 74684 27548
rect 74920 27538 74948 27911
rect 74908 27532 74960 27538
rect 74908 27474 74960 27480
rect 74540 27328 74592 27334
rect 74632 27328 74684 27334
rect 74592 27288 74632 27316
rect 74540 27270 74592 27276
rect 74632 27270 74684 27276
rect 74814 27160 74870 27169
rect 74552 27130 74764 27146
rect 74540 27124 74776 27130
rect 74592 27118 74724 27124
rect 74540 27066 74592 27072
rect 74814 27095 74870 27104
rect 74724 27066 74776 27072
rect 74828 26994 74856 27095
rect 75012 27062 75040 27950
rect 75000 27056 75052 27062
rect 75000 26998 75052 27004
rect 74448 26988 74500 26994
rect 74448 26930 74500 26936
rect 74816 26988 74868 26994
rect 74816 26930 74868 26936
rect 74570 26684 74878 26693
rect 74570 26682 74576 26684
rect 74632 26682 74656 26684
rect 74712 26682 74736 26684
rect 74792 26682 74816 26684
rect 74872 26682 74878 26684
rect 74632 26630 74634 26682
rect 74814 26630 74816 26682
rect 74570 26628 74576 26630
rect 74632 26628 74656 26630
rect 74712 26628 74736 26630
rect 74792 26628 74816 26630
rect 74872 26628 74878 26630
rect 74570 26619 74878 26628
rect 74908 26580 74960 26586
rect 74908 26522 74960 26528
rect 74724 26512 74776 26518
rect 74724 26454 74776 26460
rect 74736 26246 74764 26454
rect 74920 26382 74948 26522
rect 75104 26382 75132 29294
rect 76010 29294 76328 29322
rect 76010 29200 76066 29294
rect 75276 28076 75328 28082
rect 75276 28018 75328 28024
rect 75182 27704 75238 27713
rect 75182 27639 75238 27648
rect 75196 27538 75224 27639
rect 75288 27606 75316 28018
rect 76196 27940 76248 27946
rect 76196 27882 76248 27888
rect 75920 27872 75972 27878
rect 75920 27814 75972 27820
rect 75276 27600 75328 27606
rect 75276 27542 75328 27548
rect 75184 27532 75236 27538
rect 75184 27474 75236 27480
rect 75932 27470 75960 27814
rect 75920 27464 75972 27470
rect 75920 27406 75972 27412
rect 76012 27328 76064 27334
rect 75932 27288 76012 27316
rect 75932 26926 75960 27288
rect 76012 27270 76064 27276
rect 76208 26926 76236 27882
rect 75920 26920 75972 26926
rect 75550 26888 75606 26897
rect 75920 26862 75972 26868
rect 76104 26920 76156 26926
rect 76104 26862 76156 26868
rect 76196 26920 76248 26926
rect 76196 26862 76248 26868
rect 75550 26823 75606 26832
rect 75564 26790 75592 26823
rect 75552 26784 75604 26790
rect 75552 26726 75604 26732
rect 74908 26376 74960 26382
rect 74908 26318 74960 26324
rect 75092 26376 75144 26382
rect 75092 26318 75144 26324
rect 74724 26240 74776 26246
rect 74724 26182 74776 26188
rect 76116 26042 76144 26862
rect 76104 26036 76156 26042
rect 76104 25978 76156 25984
rect 76300 25906 76328 29294
rect 76654 29294 76788 29322
rect 76654 29200 76710 29294
rect 76760 27470 76788 29294
rect 77298 29294 77432 29322
rect 77298 29200 77354 29294
rect 76748 27464 76800 27470
rect 76748 27406 76800 27412
rect 76840 27464 76892 27470
rect 76840 27406 76892 27412
rect 76562 27160 76618 27169
rect 76562 27095 76618 27104
rect 76576 27062 76604 27095
rect 76564 27056 76616 27062
rect 76564 26998 76616 27004
rect 76472 26784 76524 26790
rect 76472 26726 76524 26732
rect 76564 26784 76616 26790
rect 76564 26726 76616 26732
rect 76484 26382 76512 26726
rect 76576 26586 76604 26726
rect 76564 26580 76616 26586
rect 76564 26522 76616 26528
rect 76472 26376 76524 26382
rect 76472 26318 76524 26324
rect 76656 26240 76708 26246
rect 76656 26182 76708 26188
rect 76288 25900 76340 25906
rect 76288 25842 76340 25848
rect 74570 25596 74878 25605
rect 74570 25594 74576 25596
rect 74632 25594 74656 25596
rect 74712 25594 74736 25596
rect 74792 25594 74816 25596
rect 74872 25594 74878 25596
rect 74632 25542 74634 25594
rect 74814 25542 74816 25594
rect 74570 25540 74576 25542
rect 74632 25540 74656 25542
rect 74712 25540 74736 25542
rect 74792 25540 74816 25542
rect 74872 25540 74878 25542
rect 74570 25531 74878 25540
rect 74570 24508 74878 24517
rect 74570 24506 74576 24508
rect 74632 24506 74656 24508
rect 74712 24506 74736 24508
rect 74792 24506 74816 24508
rect 74872 24506 74878 24508
rect 74632 24454 74634 24506
rect 74814 24454 74816 24506
rect 74570 24452 74576 24454
rect 74632 24452 74656 24454
rect 74712 24452 74736 24454
rect 74792 24452 74816 24454
rect 74872 24452 74878 24454
rect 74570 24443 74878 24452
rect 74570 23420 74878 23429
rect 74570 23418 74576 23420
rect 74632 23418 74656 23420
rect 74712 23418 74736 23420
rect 74792 23418 74816 23420
rect 74872 23418 74878 23420
rect 74632 23366 74634 23418
rect 74814 23366 74816 23418
rect 74570 23364 74576 23366
rect 74632 23364 74656 23366
rect 74712 23364 74736 23366
rect 74792 23364 74816 23366
rect 74872 23364 74878 23366
rect 74570 23355 74878 23364
rect 74570 22332 74878 22341
rect 74570 22330 74576 22332
rect 74632 22330 74656 22332
rect 74712 22330 74736 22332
rect 74792 22330 74816 22332
rect 74872 22330 74878 22332
rect 74632 22278 74634 22330
rect 74814 22278 74816 22330
rect 74570 22276 74576 22278
rect 74632 22276 74656 22278
rect 74712 22276 74736 22278
rect 74792 22276 74816 22278
rect 74872 22276 74878 22278
rect 74570 22267 74878 22276
rect 74570 21244 74878 21253
rect 74570 21242 74576 21244
rect 74632 21242 74656 21244
rect 74712 21242 74736 21244
rect 74792 21242 74816 21244
rect 74872 21242 74878 21244
rect 74632 21190 74634 21242
rect 74814 21190 74816 21242
rect 74570 21188 74576 21190
rect 74632 21188 74656 21190
rect 74712 21188 74736 21190
rect 74792 21188 74816 21190
rect 74872 21188 74878 21190
rect 74570 21179 74878 21188
rect 74570 20156 74878 20165
rect 74570 20154 74576 20156
rect 74632 20154 74656 20156
rect 74712 20154 74736 20156
rect 74792 20154 74816 20156
rect 74872 20154 74878 20156
rect 74632 20102 74634 20154
rect 74814 20102 74816 20154
rect 74570 20100 74576 20102
rect 74632 20100 74656 20102
rect 74712 20100 74736 20102
rect 74792 20100 74816 20102
rect 74872 20100 74878 20102
rect 74570 20091 74878 20100
rect 74570 19068 74878 19077
rect 74570 19066 74576 19068
rect 74632 19066 74656 19068
rect 74712 19066 74736 19068
rect 74792 19066 74816 19068
rect 74872 19066 74878 19068
rect 74632 19014 74634 19066
rect 74814 19014 74816 19066
rect 74570 19012 74576 19014
rect 74632 19012 74656 19014
rect 74712 19012 74736 19014
rect 74792 19012 74816 19014
rect 74872 19012 74878 19014
rect 74570 19003 74878 19012
rect 74570 17980 74878 17989
rect 74570 17978 74576 17980
rect 74632 17978 74656 17980
rect 74712 17978 74736 17980
rect 74792 17978 74816 17980
rect 74872 17978 74878 17980
rect 74632 17926 74634 17978
rect 74814 17926 74816 17978
rect 74570 17924 74576 17926
rect 74632 17924 74656 17926
rect 74712 17924 74736 17926
rect 74792 17924 74816 17926
rect 74872 17924 74878 17926
rect 74570 17915 74878 17924
rect 74570 16892 74878 16901
rect 74570 16890 74576 16892
rect 74632 16890 74656 16892
rect 74712 16890 74736 16892
rect 74792 16890 74816 16892
rect 74872 16890 74878 16892
rect 74632 16838 74634 16890
rect 74814 16838 74816 16890
rect 74570 16836 74576 16838
rect 74632 16836 74656 16838
rect 74712 16836 74736 16838
rect 74792 16836 74816 16838
rect 74872 16836 74878 16838
rect 74570 16827 74878 16836
rect 74570 15804 74878 15813
rect 74570 15802 74576 15804
rect 74632 15802 74656 15804
rect 74712 15802 74736 15804
rect 74792 15802 74816 15804
rect 74872 15802 74878 15804
rect 74632 15750 74634 15802
rect 74814 15750 74816 15802
rect 74570 15748 74576 15750
rect 74632 15748 74656 15750
rect 74712 15748 74736 15750
rect 74792 15748 74816 15750
rect 74872 15748 74878 15750
rect 74570 15739 74878 15748
rect 74570 14716 74878 14725
rect 74570 14714 74576 14716
rect 74632 14714 74656 14716
rect 74712 14714 74736 14716
rect 74792 14714 74816 14716
rect 74872 14714 74878 14716
rect 74632 14662 74634 14714
rect 74814 14662 74816 14714
rect 74570 14660 74576 14662
rect 74632 14660 74656 14662
rect 74712 14660 74736 14662
rect 74792 14660 74816 14662
rect 74872 14660 74878 14662
rect 74570 14651 74878 14660
rect 74570 13628 74878 13637
rect 74570 13626 74576 13628
rect 74632 13626 74656 13628
rect 74712 13626 74736 13628
rect 74792 13626 74816 13628
rect 74872 13626 74878 13628
rect 74632 13574 74634 13626
rect 74814 13574 74816 13626
rect 74570 13572 74576 13574
rect 74632 13572 74656 13574
rect 74712 13572 74736 13574
rect 74792 13572 74816 13574
rect 74872 13572 74878 13574
rect 74570 13563 74878 13572
rect 73804 12980 73856 12986
rect 73804 12922 73856 12928
rect 76380 12640 76432 12646
rect 76380 12582 76432 12588
rect 74570 12540 74878 12549
rect 74570 12538 74576 12540
rect 74632 12538 74656 12540
rect 74712 12538 74736 12540
rect 74792 12538 74816 12540
rect 74872 12538 74878 12540
rect 74632 12486 74634 12538
rect 74814 12486 74816 12538
rect 74570 12484 74576 12486
rect 74632 12484 74656 12486
rect 74712 12484 74736 12486
rect 74792 12484 74816 12486
rect 74872 12484 74878 12486
rect 74570 12475 74878 12484
rect 75552 11892 75604 11898
rect 75552 11834 75604 11840
rect 74570 11452 74878 11461
rect 74570 11450 74576 11452
rect 74632 11450 74656 11452
rect 74712 11450 74736 11452
rect 74792 11450 74816 11452
rect 74872 11450 74878 11452
rect 74632 11398 74634 11450
rect 74814 11398 74816 11450
rect 74570 11396 74576 11398
rect 74632 11396 74656 11398
rect 74712 11396 74736 11398
rect 74792 11396 74816 11398
rect 74872 11396 74878 11398
rect 74570 11387 74878 11396
rect 74570 10364 74878 10373
rect 74570 10362 74576 10364
rect 74632 10362 74656 10364
rect 74712 10362 74736 10364
rect 74792 10362 74816 10364
rect 74872 10362 74878 10364
rect 74632 10310 74634 10362
rect 74814 10310 74816 10362
rect 74570 10308 74576 10310
rect 74632 10308 74656 10310
rect 74712 10308 74736 10310
rect 74792 10308 74816 10310
rect 74872 10308 74878 10310
rect 74570 10299 74878 10308
rect 74570 9276 74878 9285
rect 74570 9274 74576 9276
rect 74632 9274 74656 9276
rect 74712 9274 74736 9276
rect 74792 9274 74816 9276
rect 74872 9274 74878 9276
rect 74632 9222 74634 9274
rect 74814 9222 74816 9274
rect 74570 9220 74576 9222
rect 74632 9220 74656 9222
rect 74712 9220 74736 9222
rect 74792 9220 74816 9222
rect 74872 9220 74878 9222
rect 74570 9211 74878 9220
rect 74570 8188 74878 8197
rect 74570 8186 74576 8188
rect 74632 8186 74656 8188
rect 74712 8186 74736 8188
rect 74792 8186 74816 8188
rect 74872 8186 74878 8188
rect 74632 8134 74634 8186
rect 74814 8134 74816 8186
rect 74570 8132 74576 8134
rect 74632 8132 74656 8134
rect 74712 8132 74736 8134
rect 74792 8132 74816 8134
rect 74872 8132 74878 8134
rect 74570 8123 74878 8132
rect 74570 7100 74878 7109
rect 74570 7098 74576 7100
rect 74632 7098 74656 7100
rect 74712 7098 74736 7100
rect 74792 7098 74816 7100
rect 74872 7098 74878 7100
rect 74632 7046 74634 7098
rect 74814 7046 74816 7098
rect 74570 7044 74576 7046
rect 74632 7044 74656 7046
rect 74712 7044 74736 7046
rect 74792 7044 74816 7046
rect 74872 7044 74878 7046
rect 74570 7035 74878 7044
rect 74570 6012 74878 6021
rect 74570 6010 74576 6012
rect 74632 6010 74656 6012
rect 74712 6010 74736 6012
rect 74792 6010 74816 6012
rect 74872 6010 74878 6012
rect 74632 5958 74634 6010
rect 74814 5958 74816 6010
rect 74570 5956 74576 5958
rect 74632 5956 74656 5958
rect 74712 5956 74736 5958
rect 74792 5956 74816 5958
rect 74872 5956 74878 5958
rect 74570 5947 74878 5956
rect 74570 4924 74878 4933
rect 74570 4922 74576 4924
rect 74632 4922 74656 4924
rect 74712 4922 74736 4924
rect 74792 4922 74816 4924
rect 74872 4922 74878 4924
rect 74632 4870 74634 4922
rect 74814 4870 74816 4922
rect 74570 4868 74576 4870
rect 74632 4868 74656 4870
rect 74712 4868 74736 4870
rect 74792 4868 74816 4870
rect 74872 4868 74878 4870
rect 74570 4859 74878 4868
rect 73068 4208 73120 4214
rect 73068 4150 73120 4156
rect 73080 3942 73108 4150
rect 74184 4010 74396 4026
rect 74172 4004 74408 4010
rect 74224 3998 74356 4004
rect 74172 3946 74224 3952
rect 74356 3946 74408 3952
rect 73068 3936 73120 3942
rect 73068 3878 73120 3884
rect 73160 3936 73212 3942
rect 73160 3878 73212 3884
rect 73712 3936 73764 3942
rect 73712 3878 73764 3884
rect 74080 3936 74132 3942
rect 74080 3878 74132 3884
rect 73068 3664 73120 3670
rect 73068 3606 73120 3612
rect 72882 1728 72938 1737
rect 72882 1663 72938 1672
rect 72804 870 72924 898
rect 72804 800 72832 870
rect 61304 734 61516 762
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 72896 762 72924 870
rect 73080 762 73108 3606
rect 73172 3534 73200 3878
rect 73160 3528 73212 3534
rect 73160 3470 73212 3476
rect 73436 2848 73488 2854
rect 73434 2816 73436 2825
rect 73488 2816 73490 2825
rect 73434 2751 73490 2760
rect 73528 2508 73580 2514
rect 73528 2450 73580 2456
rect 73540 2106 73568 2450
rect 73724 2446 73752 3878
rect 74092 3670 74120 3878
rect 74570 3836 74878 3845
rect 74570 3834 74576 3836
rect 74632 3834 74656 3836
rect 74712 3834 74736 3836
rect 74792 3834 74816 3836
rect 74872 3834 74878 3836
rect 74632 3782 74634 3834
rect 74814 3782 74816 3834
rect 74570 3780 74576 3782
rect 74632 3780 74656 3782
rect 74712 3780 74736 3782
rect 74792 3780 74816 3782
rect 74872 3780 74878 3782
rect 74570 3771 74878 3780
rect 74080 3664 74132 3670
rect 74080 3606 74132 3612
rect 74172 3528 74224 3534
rect 74172 3470 74224 3476
rect 74908 3528 74960 3534
rect 74908 3470 74960 3476
rect 74184 3398 74212 3470
rect 74172 3392 74224 3398
rect 74172 3334 74224 3340
rect 74540 3392 74592 3398
rect 74540 3334 74592 3340
rect 74552 3126 74580 3334
rect 74540 3120 74592 3126
rect 74540 3062 74592 3068
rect 74570 2748 74878 2757
rect 74570 2746 74576 2748
rect 74632 2746 74656 2748
rect 74712 2746 74736 2748
rect 74792 2746 74816 2748
rect 74872 2746 74878 2748
rect 74632 2694 74634 2746
rect 74814 2694 74816 2746
rect 74570 2692 74576 2694
rect 74632 2692 74656 2694
rect 74712 2692 74736 2694
rect 74792 2692 74816 2694
rect 74872 2692 74878 2694
rect 74570 2683 74878 2692
rect 74630 2544 74686 2553
rect 73988 2508 74040 2514
rect 73908 2468 73988 2496
rect 73712 2440 73764 2446
rect 73712 2382 73764 2388
rect 73620 2304 73672 2310
rect 73620 2246 73672 2252
rect 73632 2106 73660 2246
rect 73528 2100 73580 2106
rect 73528 2042 73580 2048
rect 73620 2100 73672 2106
rect 73620 2042 73672 2048
rect 73908 1970 73936 2468
rect 74630 2479 74686 2488
rect 73988 2450 74040 2456
rect 74644 2310 74672 2479
rect 74632 2304 74684 2310
rect 74632 2246 74684 2252
rect 73896 1964 73948 1970
rect 73896 1906 73948 1912
rect 73988 1964 74040 1970
rect 73988 1906 74040 1912
rect 74000 1698 74028 1906
rect 73988 1692 74040 1698
rect 73988 1634 74040 1640
rect 74080 1692 74132 1698
rect 74080 1634 74132 1640
rect 74092 800 74120 1634
rect 74920 1442 74948 3470
rect 75460 3392 75512 3398
rect 75460 3334 75512 3340
rect 75368 3120 75420 3126
rect 75368 3062 75420 3068
rect 75092 2916 75144 2922
rect 75092 2858 75144 2864
rect 75104 1698 75132 2858
rect 75380 1902 75408 3062
rect 75368 1896 75420 1902
rect 75368 1838 75420 1844
rect 75092 1692 75144 1698
rect 75092 1634 75144 1640
rect 74736 1414 74948 1442
rect 74736 800 74764 1414
rect 75472 1034 75500 3334
rect 75564 2854 75592 11834
rect 76392 11830 76420 12582
rect 76380 11824 76432 11830
rect 76380 11766 76432 11772
rect 76668 8974 76696 26182
rect 76852 25838 76880 27406
rect 77300 27124 77352 27130
rect 77300 27066 77352 27072
rect 76840 25832 76892 25838
rect 76840 25774 76892 25780
rect 77312 22094 77340 27066
rect 77404 26586 77432 29294
rect 78586 29200 78642 30000
rect 79230 29200 79286 30000
rect 80518 29200 80574 30000
rect 81162 29322 81218 30000
rect 82450 29322 82506 30000
rect 83094 29322 83150 30000
rect 83738 29322 83794 30000
rect 85026 29322 85082 30000
rect 81162 29294 81388 29322
rect 81162 29200 81218 29294
rect 78600 27878 78628 29200
rect 78588 27872 78640 27878
rect 78588 27814 78640 27820
rect 78864 27532 78916 27538
rect 78864 27474 78916 27480
rect 78772 27396 78824 27402
rect 78772 27338 78824 27344
rect 78588 27328 78640 27334
rect 78586 27296 78588 27305
rect 78640 27296 78642 27305
rect 78586 27231 78642 27240
rect 78680 26852 78732 26858
rect 78680 26794 78732 26800
rect 78404 26784 78456 26790
rect 78404 26726 78456 26732
rect 78416 26586 78444 26726
rect 77392 26580 77444 26586
rect 77392 26522 77444 26528
rect 78404 26580 78456 26586
rect 78404 26522 78456 26528
rect 77484 26444 77536 26450
rect 77484 26386 77536 26392
rect 77496 26042 77524 26386
rect 78692 26382 78720 26794
rect 78784 26625 78812 27338
rect 78770 26616 78826 26625
rect 78770 26551 78826 26560
rect 77576 26376 77628 26382
rect 77576 26318 77628 26324
rect 78680 26376 78732 26382
rect 78680 26318 78732 26324
rect 77484 26036 77536 26042
rect 77484 25978 77536 25984
rect 77588 25906 77616 26318
rect 77576 25900 77628 25906
rect 77576 25842 77628 25848
rect 78876 25702 78904 27474
rect 79046 27432 79102 27441
rect 79046 27367 79102 27376
rect 79060 27334 79088 27367
rect 78956 27328 79008 27334
rect 78956 27270 79008 27276
rect 79048 27328 79100 27334
rect 79048 27270 79100 27276
rect 78864 25696 78916 25702
rect 78864 25638 78916 25644
rect 77312 22066 77524 22094
rect 77024 12776 77076 12782
rect 77024 12718 77076 12724
rect 77036 11694 77064 12718
rect 77024 11688 77076 11694
rect 77024 11630 77076 11636
rect 76656 8968 76708 8974
rect 76656 8910 76708 8916
rect 76472 7812 76524 7818
rect 76472 7754 76524 7760
rect 76012 3392 76064 3398
rect 76012 3334 76064 3340
rect 76024 3194 76052 3334
rect 76012 3188 76064 3194
rect 76012 3130 76064 3136
rect 76484 2922 76512 7754
rect 77036 4162 77064 11630
rect 77208 8492 77260 8498
rect 77208 8434 77260 8440
rect 77220 8022 77248 8434
rect 77208 8016 77260 8022
rect 77208 7958 77260 7964
rect 76944 4134 77064 4162
rect 77208 4140 77260 4146
rect 76840 3052 76892 3058
rect 76840 2994 76892 3000
rect 76852 2922 76880 2994
rect 76944 2990 76972 4134
rect 77208 4082 77260 4088
rect 77024 3936 77076 3942
rect 77024 3878 77076 3884
rect 77036 3126 77064 3878
rect 77116 3392 77168 3398
rect 77116 3334 77168 3340
rect 77128 3194 77156 3334
rect 77116 3188 77168 3194
rect 77116 3130 77168 3136
rect 77024 3120 77076 3126
rect 77024 3062 77076 3068
rect 77114 3088 77170 3097
rect 77114 3023 77170 3032
rect 77128 2990 77156 3023
rect 76932 2984 76984 2990
rect 76932 2926 76984 2932
rect 77116 2984 77168 2990
rect 77116 2926 77168 2932
rect 75736 2916 75788 2922
rect 75736 2858 75788 2864
rect 76472 2916 76524 2922
rect 76472 2858 76524 2864
rect 76840 2916 76892 2922
rect 76840 2858 76892 2864
rect 75552 2848 75604 2854
rect 75552 2790 75604 2796
rect 75748 2428 75776 2858
rect 76944 2774 76972 2926
rect 77220 2825 77248 4082
rect 77496 3398 77524 22066
rect 78036 20324 78088 20330
rect 78036 20266 78088 20272
rect 78048 3534 78076 20266
rect 78680 20256 78732 20262
rect 78680 20198 78732 20204
rect 78692 19854 78720 20198
rect 78680 19848 78732 19854
rect 78680 19790 78732 19796
rect 78968 19786 78996 27270
rect 79244 27130 79272 29200
rect 79600 27872 79652 27878
rect 79600 27814 79652 27820
rect 79784 27872 79836 27878
rect 79784 27814 79836 27820
rect 80428 27872 80480 27878
rect 80428 27814 80480 27820
rect 79414 27704 79470 27713
rect 79414 27639 79470 27648
rect 79428 27538 79456 27639
rect 79416 27532 79468 27538
rect 79416 27474 79468 27480
rect 79324 27328 79376 27334
rect 79324 27270 79376 27276
rect 79336 27169 79364 27270
rect 79322 27160 79378 27169
rect 79232 27124 79284 27130
rect 79322 27095 79378 27104
rect 79232 27066 79284 27072
rect 79428 27044 79456 27474
rect 79612 27470 79640 27814
rect 79796 27606 79824 27814
rect 79784 27600 79836 27606
rect 79784 27542 79836 27548
rect 79600 27464 79652 27470
rect 79600 27406 79652 27412
rect 80242 27296 80298 27305
rect 80242 27231 80298 27240
rect 79876 27124 79928 27130
rect 79876 27066 79928 27072
rect 79336 27016 79456 27044
rect 79048 26988 79100 26994
rect 79048 26930 79100 26936
rect 79060 26518 79088 26930
rect 79336 26772 79364 27016
rect 79244 26744 79364 26772
rect 79508 26784 79560 26790
rect 79048 26512 79100 26518
rect 79048 26454 79100 26460
rect 79244 21486 79272 26744
rect 79508 26726 79560 26732
rect 79520 26586 79548 26726
rect 79888 26602 79916 27066
rect 80060 26988 80112 26994
rect 80060 26930 80112 26936
rect 80072 26897 80100 26930
rect 80256 26897 80284 27231
rect 80334 27160 80390 27169
rect 80334 27095 80390 27104
rect 80058 26888 80114 26897
rect 80058 26823 80114 26832
rect 80242 26888 80298 26897
rect 80242 26823 80298 26832
rect 79508 26580 79560 26586
rect 79508 26522 79560 26528
rect 79796 26574 79916 26602
rect 79690 26480 79746 26489
rect 79690 26415 79746 26424
rect 79704 26382 79732 26415
rect 79692 26376 79744 26382
rect 79692 26318 79744 26324
rect 79600 26240 79652 26246
rect 79796 26217 79824 26574
rect 80242 26344 80298 26353
rect 80348 26330 80376 27095
rect 80440 26353 80468 27814
rect 80532 27470 80560 29200
rect 81256 27600 81308 27606
rect 81176 27560 81256 27588
rect 80520 27464 80572 27470
rect 80520 27406 80572 27412
rect 81176 26761 81204 27560
rect 81360 27588 81388 29294
rect 82450 29294 82584 29322
rect 82450 29200 82506 29294
rect 82556 27606 82584 29294
rect 83094 29294 83688 29322
rect 83094 29200 83150 29294
rect 81440 27600 81492 27606
rect 81360 27560 81440 27588
rect 81256 27542 81308 27548
rect 81440 27542 81492 27548
rect 82544 27600 82596 27606
rect 82544 27542 82596 27548
rect 81992 27464 82044 27470
rect 81992 27406 82044 27412
rect 82728 27464 82780 27470
rect 83660 27452 83688 29294
rect 83738 29294 84056 29322
rect 83738 29200 83794 29294
rect 83740 27464 83792 27470
rect 83660 27424 83740 27452
rect 82728 27406 82780 27412
rect 83740 27406 83792 27412
rect 83924 27464 83976 27470
rect 83924 27406 83976 27412
rect 81162 26752 81218 26761
rect 81162 26687 81218 26696
rect 81898 26616 81954 26625
rect 81898 26551 81954 26560
rect 81438 26480 81494 26489
rect 81438 26415 81494 26424
rect 80298 26302 80376 26330
rect 80426 26344 80482 26353
rect 80242 26279 80298 26288
rect 80426 26279 80482 26288
rect 81164 26308 81216 26314
rect 81164 26250 81216 26256
rect 79600 26182 79652 26188
rect 79782 26208 79838 26217
rect 79232 21480 79284 21486
rect 79232 21422 79284 21428
rect 79048 20460 79100 20466
rect 79048 20402 79100 20408
rect 79060 20058 79088 20402
rect 79244 20398 79272 21422
rect 79232 20392 79284 20398
rect 79232 20334 79284 20340
rect 79048 20052 79100 20058
rect 79048 19994 79100 20000
rect 78956 19780 79008 19786
rect 78956 19722 79008 19728
rect 79232 4616 79284 4622
rect 79232 4558 79284 4564
rect 79244 4146 79272 4558
rect 79232 4140 79284 4146
rect 79232 4082 79284 4088
rect 79508 3936 79560 3942
rect 79508 3878 79560 3884
rect 78036 3528 78088 3534
rect 78036 3470 78088 3476
rect 77484 3392 77536 3398
rect 77484 3334 77536 3340
rect 77300 3052 77352 3058
rect 77300 2994 77352 3000
rect 77206 2816 77262 2825
rect 76944 2746 77064 2774
rect 77206 2751 77262 2760
rect 77036 2514 77064 2746
rect 77024 2508 77076 2514
rect 77024 2450 77076 2456
rect 77208 2508 77260 2514
rect 77208 2450 77260 2456
rect 75828 2440 75880 2446
rect 75748 2400 75828 2428
rect 75828 2382 75880 2388
rect 76840 2304 76892 2310
rect 76840 2246 76892 2252
rect 77116 2304 77168 2310
rect 77116 2246 77168 2252
rect 75552 1896 75604 1902
rect 75550 1864 75552 1873
rect 75604 1864 75606 1873
rect 75550 1799 75606 1808
rect 76852 1766 76880 2246
rect 76840 1760 76892 1766
rect 76840 1702 76892 1708
rect 75380 1006 75500 1034
rect 75380 800 75408 1006
rect 76668 870 76788 898
rect 76668 800 76696 870
rect 72896 734 73108 762
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 76760 762 76788 870
rect 77128 762 77156 2246
rect 77220 1902 77248 2450
rect 77208 1896 77260 1902
rect 77208 1838 77260 1844
rect 77312 800 77340 2994
rect 78034 2816 78090 2825
rect 78034 2751 78090 2760
rect 78048 2446 78076 2751
rect 79520 2446 79548 3878
rect 77392 2440 77444 2446
rect 77392 2382 77444 2388
rect 78036 2440 78088 2446
rect 78036 2382 78088 2388
rect 79508 2440 79560 2446
rect 79508 2382 79560 2388
rect 77404 2310 77432 2382
rect 77392 2304 77444 2310
rect 77392 2246 77444 2252
rect 77760 2304 77812 2310
rect 77760 2246 77812 2252
rect 78588 2304 78640 2310
rect 78588 2246 78640 2252
rect 79232 2304 79284 2310
rect 79612 2281 79640 26182
rect 79782 26143 79838 26152
rect 81176 25974 81204 26250
rect 81164 25968 81216 25974
rect 81164 25910 81216 25916
rect 80704 19712 80756 19718
rect 80704 19654 80756 19660
rect 80716 3058 80744 19654
rect 81452 17814 81480 26415
rect 81912 26382 81940 26551
rect 81900 26376 81952 26382
rect 81900 26318 81952 26324
rect 81440 17808 81492 17814
rect 81440 17750 81492 17756
rect 82004 13870 82032 27406
rect 82268 26444 82320 26450
rect 82268 26386 82320 26392
rect 82280 25906 82308 26386
rect 82268 25900 82320 25906
rect 82268 25842 82320 25848
rect 82740 21418 82768 27406
rect 83936 27130 83964 27406
rect 83924 27124 83976 27130
rect 84028 27112 84056 29294
rect 85026 29294 85528 29322
rect 85026 29200 85082 29294
rect 85210 27976 85266 27985
rect 85210 27911 85266 27920
rect 84844 27872 84896 27878
rect 84844 27814 84896 27820
rect 84856 27674 84884 27814
rect 84844 27668 84896 27674
rect 84844 27610 84896 27616
rect 85224 27538 85252 27911
rect 85500 27588 85528 29294
rect 85670 29200 85726 30000
rect 86958 29322 87014 30000
rect 87602 29322 87658 30000
rect 86958 29294 87092 29322
rect 86958 29200 87014 29294
rect 85580 27600 85632 27606
rect 85500 27560 85580 27588
rect 85580 27542 85632 27548
rect 84292 27532 84344 27538
rect 84292 27474 84344 27480
rect 85028 27532 85080 27538
rect 85028 27474 85080 27480
rect 85212 27532 85264 27538
rect 85212 27474 85264 27480
rect 84304 27334 84332 27474
rect 84292 27328 84344 27334
rect 84476 27328 84528 27334
rect 84292 27270 84344 27276
rect 84474 27296 84476 27305
rect 84528 27296 84530 27305
rect 84474 27231 84530 27240
rect 84200 27124 84252 27130
rect 84028 27084 84200 27112
rect 83924 27066 83976 27072
rect 84200 27066 84252 27072
rect 84936 27124 84988 27130
rect 84936 27066 84988 27072
rect 84016 26988 84068 26994
rect 84016 26930 84068 26936
rect 84028 26586 84056 26930
rect 84844 26920 84896 26926
rect 84948 26908 84976 27066
rect 84896 26880 84976 26908
rect 84844 26862 84896 26868
rect 84568 26852 84620 26858
rect 84568 26794 84620 26800
rect 84016 26580 84068 26586
rect 84016 26522 84068 26528
rect 82728 21412 82780 21418
rect 82728 21354 82780 21360
rect 84476 20800 84528 20806
rect 84476 20742 84528 20748
rect 84488 20466 84516 20742
rect 84476 20460 84528 20466
rect 84476 20402 84528 20408
rect 82728 17808 82780 17814
rect 82728 17750 82780 17756
rect 82740 16658 82768 17750
rect 82912 17196 82964 17202
rect 82912 17138 82964 17144
rect 82728 16652 82780 16658
rect 82728 16594 82780 16600
rect 81992 13864 82044 13870
rect 81992 13806 82044 13812
rect 82544 10736 82596 10742
rect 82544 10678 82596 10684
rect 80704 3052 80756 3058
rect 80704 2994 80756 3000
rect 81164 2848 81216 2854
rect 81164 2790 81216 2796
rect 80520 2440 80572 2446
rect 80520 2382 80572 2388
rect 79232 2246 79284 2252
rect 79598 2272 79654 2281
rect 77390 2000 77446 2009
rect 77390 1935 77446 1944
rect 77404 1902 77432 1935
rect 77392 1896 77444 1902
rect 77392 1838 77444 1844
rect 77772 1698 77800 2246
rect 77850 1728 77906 1737
rect 77760 1692 77812 1698
rect 77850 1663 77852 1672
rect 77760 1634 77812 1640
rect 77904 1663 77906 1672
rect 77852 1634 77904 1640
rect 78600 800 78628 2246
rect 79244 800 79272 2246
rect 79598 2207 79654 2216
rect 80150 2272 80206 2281
rect 80150 2207 80206 2216
rect 80058 1456 80114 1465
rect 80164 1426 80192 2207
rect 80058 1391 80060 1400
rect 80112 1391 80114 1400
rect 80152 1420 80204 1426
rect 80060 1362 80112 1368
rect 80152 1362 80204 1368
rect 80532 800 80560 2382
rect 81176 800 81204 2790
rect 82556 2650 82584 10678
rect 82636 4276 82688 4282
rect 82636 4218 82688 4224
rect 82648 4010 82676 4218
rect 82740 4078 82768 16594
rect 82924 16454 82952 17138
rect 82912 16448 82964 16454
rect 82912 16390 82964 16396
rect 83004 10464 83056 10470
rect 83004 10406 83056 10412
rect 83016 5302 83044 10406
rect 83004 5296 83056 5302
rect 83004 5238 83056 5244
rect 82820 5228 82872 5234
rect 82820 5170 82872 5176
rect 82728 4072 82780 4078
rect 82728 4014 82780 4020
rect 82636 4004 82688 4010
rect 82636 3946 82688 3952
rect 82832 3942 82860 5170
rect 82820 3936 82872 3942
rect 82820 3878 82872 3884
rect 82452 2644 82504 2650
rect 82452 2586 82504 2592
rect 82544 2644 82596 2650
rect 82728 2644 82780 2650
rect 82544 2586 82596 2592
rect 82648 2604 82728 2632
rect 82464 2530 82492 2586
rect 82648 2530 82676 2604
rect 82728 2586 82780 2592
rect 81544 2502 82124 2530
rect 82464 2502 82676 2530
rect 81348 2440 81400 2446
rect 81348 2382 81400 2388
rect 81360 1222 81388 2382
rect 81544 2378 81572 2502
rect 81992 2440 82044 2446
rect 81992 2382 82044 2388
rect 81532 2372 81584 2378
rect 81532 2314 81584 2320
rect 82004 1306 82032 2382
rect 82096 2378 82124 2502
rect 84580 2446 84608 26794
rect 85040 26042 85068 27474
rect 85210 27296 85266 27305
rect 85210 27231 85266 27240
rect 85224 26926 85252 27231
rect 85684 27062 85712 29200
rect 87064 27606 87092 29294
rect 87602 29294 87736 29322
rect 87602 29200 87658 29294
rect 87708 27606 87736 29294
rect 88246 29200 88302 30000
rect 89534 29322 89590 30000
rect 90178 29322 90234 30000
rect 89534 29294 89668 29322
rect 89534 29200 89590 29294
rect 87052 27600 87104 27606
rect 87052 27542 87104 27548
rect 87696 27600 87748 27606
rect 87696 27542 87748 27548
rect 86408 27464 86460 27470
rect 86408 27406 86460 27412
rect 87236 27464 87288 27470
rect 87236 27406 87288 27412
rect 87328 27464 87380 27470
rect 88260 27452 88288 29200
rect 88340 27464 88392 27470
rect 88260 27424 88340 27452
rect 87328 27406 87380 27412
rect 88340 27406 88392 27412
rect 89074 27432 89130 27441
rect 86132 27396 86184 27402
rect 86132 27338 86184 27344
rect 85672 27056 85724 27062
rect 85672 26998 85724 27004
rect 85304 26988 85356 26994
rect 85304 26930 85356 26936
rect 85212 26920 85264 26926
rect 85212 26862 85264 26868
rect 85316 26586 85344 26930
rect 86144 26858 86172 27338
rect 86132 26852 86184 26858
rect 86132 26794 86184 26800
rect 85396 26784 85448 26790
rect 85396 26726 85448 26732
rect 86224 26784 86276 26790
rect 86224 26726 86276 26732
rect 85408 26586 85436 26726
rect 85304 26580 85356 26586
rect 85304 26522 85356 26528
rect 85396 26580 85448 26586
rect 85396 26522 85448 26528
rect 85028 26036 85080 26042
rect 85028 25978 85080 25984
rect 85040 21010 85068 25978
rect 85028 21004 85080 21010
rect 85028 20946 85080 20952
rect 86236 14074 86264 26726
rect 86420 25158 86448 27406
rect 86960 27396 87012 27402
rect 86960 27338 87012 27344
rect 86972 27062 87000 27338
rect 86960 27056 87012 27062
rect 86960 26998 87012 27004
rect 86868 26784 86920 26790
rect 86868 26726 86920 26732
rect 86408 25152 86460 25158
rect 86408 25094 86460 25100
rect 86880 20602 86908 26726
rect 86868 20596 86920 20602
rect 86868 20538 86920 20544
rect 86224 14068 86276 14074
rect 86224 14010 86276 14016
rect 86408 14000 86460 14006
rect 86408 13942 86460 13948
rect 86420 13870 86448 13942
rect 86316 13864 86368 13870
rect 86316 13806 86368 13812
rect 86408 13864 86460 13870
rect 86408 13806 86460 13812
rect 85488 4208 85540 4214
rect 85488 4150 85540 4156
rect 85304 3188 85356 3194
rect 85304 3130 85356 3136
rect 85316 2446 85344 3130
rect 83096 2440 83148 2446
rect 83096 2382 83148 2388
rect 84568 2440 84620 2446
rect 84568 2382 84620 2388
rect 85304 2440 85356 2446
rect 85304 2382 85356 2388
rect 82084 2372 82136 2378
rect 82084 2314 82136 2320
rect 81820 1278 82032 1306
rect 81348 1216 81400 1222
rect 81348 1158 81400 1164
rect 81820 800 81848 1278
rect 83108 800 83136 2382
rect 85500 2310 85528 4150
rect 86328 2514 86356 13806
rect 86776 13728 86828 13734
rect 86776 13670 86828 13676
rect 86788 13326 86816 13670
rect 86776 13320 86828 13326
rect 86776 13262 86828 13268
rect 86592 13184 86644 13190
rect 86592 13126 86644 13132
rect 86316 2508 86368 2514
rect 86316 2450 86368 2456
rect 85672 2440 85724 2446
rect 85672 2382 85724 2388
rect 84016 2304 84068 2310
rect 84016 2246 84068 2252
rect 85028 2304 85080 2310
rect 85028 2246 85080 2252
rect 85488 2304 85540 2310
rect 85488 2246 85540 2252
rect 83752 870 83872 898
rect 83752 800 83780 870
rect 76760 734 77156 762
rect 77298 0 77354 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 83844 762 83872 870
rect 84028 762 84056 2246
rect 85040 800 85068 2246
rect 85684 800 85712 2382
rect 86604 1426 86632 13126
rect 87248 12102 87276 27406
rect 87340 27169 87368 27406
rect 89444 27396 89496 27402
rect 89074 27367 89130 27376
rect 88800 27328 88852 27334
rect 88800 27270 88852 27276
rect 87326 27160 87382 27169
rect 87326 27095 87382 27104
rect 88812 22710 88840 27270
rect 89088 27130 89116 27367
rect 89180 27356 89444 27384
rect 89076 27124 89128 27130
rect 89076 27066 89128 27072
rect 89180 26994 89208 27356
rect 89444 27338 89496 27344
rect 89294 27228 89602 27237
rect 89294 27226 89300 27228
rect 89356 27226 89380 27228
rect 89436 27226 89460 27228
rect 89516 27226 89540 27228
rect 89596 27226 89602 27228
rect 89356 27174 89358 27226
rect 89538 27174 89540 27226
rect 89294 27172 89300 27174
rect 89356 27172 89380 27174
rect 89436 27172 89460 27174
rect 89516 27172 89540 27174
rect 89596 27172 89602 27174
rect 89294 27163 89602 27172
rect 89640 26994 89668 29294
rect 90178 29294 90312 29322
rect 90178 29200 90234 29294
rect 89720 27668 89772 27674
rect 89720 27610 89772 27616
rect 89732 27402 89760 27610
rect 89720 27396 89772 27402
rect 89720 27338 89772 27344
rect 90088 27328 90140 27334
rect 90088 27270 90140 27276
rect 90180 27328 90232 27334
rect 90180 27270 90232 27276
rect 90100 27062 90128 27270
rect 90088 27056 90140 27062
rect 90088 26998 90140 27004
rect 90192 26994 90220 27270
rect 89168 26988 89220 26994
rect 89168 26930 89220 26936
rect 89628 26988 89680 26994
rect 89628 26930 89680 26936
rect 90180 26988 90232 26994
rect 90180 26930 90232 26936
rect 90088 26784 90140 26790
rect 90088 26726 90140 26732
rect 90100 26518 90128 26726
rect 90088 26512 90140 26518
rect 89074 26480 89130 26489
rect 90088 26454 90140 26460
rect 89074 26415 89130 26424
rect 90180 26444 90232 26450
rect 89088 26382 89116 26415
rect 90180 26386 90232 26392
rect 89076 26376 89128 26382
rect 89996 26376 90048 26382
rect 89076 26318 89128 26324
rect 89180 26314 89392 26330
rect 90192 26330 90220 26386
rect 90048 26324 90220 26330
rect 89996 26318 90220 26324
rect 89168 26308 89404 26314
rect 89220 26302 89352 26308
rect 89168 26250 89220 26256
rect 90008 26302 90220 26318
rect 89352 26250 89404 26256
rect 90284 26246 90312 29294
rect 91466 29200 91522 30000
rect 92110 29322 92166 30000
rect 93398 29322 93454 30000
rect 92110 29294 92428 29322
rect 92110 29200 92166 29294
rect 90640 27532 90692 27538
rect 90640 27474 90692 27480
rect 91376 27532 91428 27538
rect 91376 27474 91428 27480
rect 90362 27160 90418 27169
rect 90362 27095 90418 27104
rect 90376 26994 90404 27095
rect 90652 26994 90680 27474
rect 91008 27328 91060 27334
rect 91008 27270 91060 27276
rect 90732 27124 90784 27130
rect 90732 27066 90784 27072
rect 90364 26988 90416 26994
rect 90364 26930 90416 26936
rect 90640 26988 90692 26994
rect 90640 26930 90692 26936
rect 90456 26376 90508 26382
rect 90456 26318 90508 26324
rect 90272 26240 90324 26246
rect 90272 26182 90324 26188
rect 89294 26140 89602 26149
rect 89294 26138 89300 26140
rect 89356 26138 89380 26140
rect 89436 26138 89460 26140
rect 89516 26138 89540 26140
rect 89596 26138 89602 26140
rect 89356 26086 89358 26138
rect 89538 26086 89540 26138
rect 89294 26084 89300 26086
rect 89356 26084 89380 26086
rect 89436 26084 89460 26086
rect 89516 26084 89540 26086
rect 89596 26084 89602 26086
rect 89294 26075 89602 26084
rect 89294 25052 89602 25061
rect 89294 25050 89300 25052
rect 89356 25050 89380 25052
rect 89436 25050 89460 25052
rect 89516 25050 89540 25052
rect 89596 25050 89602 25052
rect 89356 24998 89358 25050
rect 89538 24998 89540 25050
rect 89294 24996 89300 24998
rect 89356 24996 89380 24998
rect 89436 24996 89460 24998
rect 89516 24996 89540 24998
rect 89596 24996 89602 24998
rect 89294 24987 89602 24996
rect 89294 23964 89602 23973
rect 89294 23962 89300 23964
rect 89356 23962 89380 23964
rect 89436 23962 89460 23964
rect 89516 23962 89540 23964
rect 89596 23962 89602 23964
rect 89356 23910 89358 23962
rect 89538 23910 89540 23962
rect 89294 23908 89300 23910
rect 89356 23908 89380 23910
rect 89436 23908 89460 23910
rect 89516 23908 89540 23910
rect 89596 23908 89602 23910
rect 89294 23899 89602 23908
rect 89294 22876 89602 22885
rect 89294 22874 89300 22876
rect 89356 22874 89380 22876
rect 89436 22874 89460 22876
rect 89516 22874 89540 22876
rect 89596 22874 89602 22876
rect 89356 22822 89358 22874
rect 89538 22822 89540 22874
rect 89294 22820 89300 22822
rect 89356 22820 89380 22822
rect 89436 22820 89460 22822
rect 89516 22820 89540 22822
rect 89596 22820 89602 22822
rect 89294 22811 89602 22820
rect 88800 22704 88852 22710
rect 88800 22646 88852 22652
rect 90468 22094 90496 26318
rect 90376 22066 90496 22094
rect 89294 21788 89602 21797
rect 89294 21786 89300 21788
rect 89356 21786 89380 21788
rect 89436 21786 89460 21788
rect 89516 21786 89540 21788
rect 89596 21786 89602 21788
rect 89356 21734 89358 21786
rect 89538 21734 89540 21786
rect 89294 21732 89300 21734
rect 89356 21732 89380 21734
rect 89436 21732 89460 21734
rect 89516 21732 89540 21734
rect 89596 21732 89602 21734
rect 89294 21723 89602 21732
rect 89294 20700 89602 20709
rect 89294 20698 89300 20700
rect 89356 20698 89380 20700
rect 89436 20698 89460 20700
rect 89516 20698 89540 20700
rect 89596 20698 89602 20700
rect 89356 20646 89358 20698
rect 89538 20646 89540 20698
rect 89294 20644 89300 20646
rect 89356 20644 89380 20646
rect 89436 20644 89460 20646
rect 89516 20644 89540 20646
rect 89596 20644 89602 20646
rect 89294 20635 89602 20644
rect 89294 19612 89602 19621
rect 89294 19610 89300 19612
rect 89356 19610 89380 19612
rect 89436 19610 89460 19612
rect 89516 19610 89540 19612
rect 89596 19610 89602 19612
rect 89356 19558 89358 19610
rect 89538 19558 89540 19610
rect 89294 19556 89300 19558
rect 89356 19556 89380 19558
rect 89436 19556 89460 19558
rect 89516 19556 89540 19558
rect 89596 19556 89602 19558
rect 89294 19547 89602 19556
rect 89294 18524 89602 18533
rect 89294 18522 89300 18524
rect 89356 18522 89380 18524
rect 89436 18522 89460 18524
rect 89516 18522 89540 18524
rect 89596 18522 89602 18524
rect 89356 18470 89358 18522
rect 89538 18470 89540 18522
rect 89294 18468 89300 18470
rect 89356 18468 89380 18470
rect 89436 18468 89460 18470
rect 89516 18468 89540 18470
rect 89596 18468 89602 18470
rect 89294 18459 89602 18468
rect 89294 17436 89602 17445
rect 89294 17434 89300 17436
rect 89356 17434 89380 17436
rect 89436 17434 89460 17436
rect 89516 17434 89540 17436
rect 89596 17434 89602 17436
rect 89356 17382 89358 17434
rect 89538 17382 89540 17434
rect 89294 17380 89300 17382
rect 89356 17380 89380 17382
rect 89436 17380 89460 17382
rect 89516 17380 89540 17382
rect 89596 17380 89602 17382
rect 89294 17371 89602 17380
rect 90376 16998 90404 22066
rect 90364 16992 90416 16998
rect 90364 16934 90416 16940
rect 89294 16348 89602 16357
rect 89294 16346 89300 16348
rect 89356 16346 89380 16348
rect 89436 16346 89460 16348
rect 89516 16346 89540 16348
rect 89596 16346 89602 16348
rect 89356 16294 89358 16346
rect 89538 16294 89540 16346
rect 89294 16292 89300 16294
rect 89356 16292 89380 16294
rect 89436 16292 89460 16294
rect 89516 16292 89540 16294
rect 89596 16292 89602 16294
rect 89294 16283 89602 16292
rect 89294 15260 89602 15269
rect 89294 15258 89300 15260
rect 89356 15258 89380 15260
rect 89436 15258 89460 15260
rect 89516 15258 89540 15260
rect 89596 15258 89602 15260
rect 89356 15206 89358 15258
rect 89538 15206 89540 15258
rect 89294 15204 89300 15206
rect 89356 15204 89380 15206
rect 89436 15204 89460 15206
rect 89516 15204 89540 15206
rect 89596 15204 89602 15206
rect 89294 15195 89602 15204
rect 90652 14346 90680 26930
rect 90744 26790 90772 27066
rect 90732 26784 90784 26790
rect 90732 26726 90784 26732
rect 90916 26784 90968 26790
rect 90916 26726 90968 26732
rect 90640 14340 90692 14346
rect 90640 14282 90692 14288
rect 89294 14172 89602 14181
rect 89294 14170 89300 14172
rect 89356 14170 89380 14172
rect 89436 14170 89460 14172
rect 89516 14170 89540 14172
rect 89596 14170 89602 14172
rect 89356 14118 89358 14170
rect 89538 14118 89540 14170
rect 89294 14116 89300 14118
rect 89356 14116 89380 14118
rect 89436 14116 89460 14118
rect 89516 14116 89540 14118
rect 89596 14116 89602 14118
rect 89294 14107 89602 14116
rect 89294 13084 89602 13093
rect 89294 13082 89300 13084
rect 89356 13082 89380 13084
rect 89436 13082 89460 13084
rect 89516 13082 89540 13084
rect 89596 13082 89602 13084
rect 89356 13030 89358 13082
rect 89538 13030 89540 13082
rect 89294 13028 89300 13030
rect 89356 13028 89380 13030
rect 89436 13028 89460 13030
rect 89516 13028 89540 13030
rect 89596 13028 89602 13030
rect 89294 13019 89602 13028
rect 87236 12096 87288 12102
rect 87236 12038 87288 12044
rect 89294 11996 89602 12005
rect 89294 11994 89300 11996
rect 89356 11994 89380 11996
rect 89436 11994 89460 11996
rect 89516 11994 89540 11996
rect 89596 11994 89602 11996
rect 89356 11942 89358 11994
rect 89538 11942 89540 11994
rect 89294 11940 89300 11942
rect 89356 11940 89380 11942
rect 89436 11940 89460 11942
rect 89516 11940 89540 11942
rect 89596 11940 89602 11942
rect 89294 11931 89602 11940
rect 89294 10908 89602 10917
rect 89294 10906 89300 10908
rect 89356 10906 89380 10908
rect 89436 10906 89460 10908
rect 89516 10906 89540 10908
rect 89596 10906 89602 10908
rect 89356 10854 89358 10906
rect 89538 10854 89540 10906
rect 89294 10852 89300 10854
rect 89356 10852 89380 10854
rect 89436 10852 89460 10854
rect 89516 10852 89540 10854
rect 89596 10852 89602 10854
rect 89294 10843 89602 10852
rect 89294 9820 89602 9829
rect 89294 9818 89300 9820
rect 89356 9818 89380 9820
rect 89436 9818 89460 9820
rect 89516 9818 89540 9820
rect 89596 9818 89602 9820
rect 89356 9766 89358 9818
rect 89538 9766 89540 9818
rect 89294 9764 89300 9766
rect 89356 9764 89380 9766
rect 89436 9764 89460 9766
rect 89516 9764 89540 9766
rect 89596 9764 89602 9766
rect 89294 9755 89602 9764
rect 89294 8732 89602 8741
rect 89294 8730 89300 8732
rect 89356 8730 89380 8732
rect 89436 8730 89460 8732
rect 89516 8730 89540 8732
rect 89596 8730 89602 8732
rect 89356 8678 89358 8730
rect 89538 8678 89540 8730
rect 89294 8676 89300 8678
rect 89356 8676 89380 8678
rect 89436 8676 89460 8678
rect 89516 8676 89540 8678
rect 89596 8676 89602 8678
rect 89294 8667 89602 8676
rect 89294 7644 89602 7653
rect 89294 7642 89300 7644
rect 89356 7642 89380 7644
rect 89436 7642 89460 7644
rect 89516 7642 89540 7644
rect 89596 7642 89602 7644
rect 89356 7590 89358 7642
rect 89538 7590 89540 7642
rect 89294 7588 89300 7590
rect 89356 7588 89380 7590
rect 89436 7588 89460 7590
rect 89516 7588 89540 7590
rect 89596 7588 89602 7590
rect 89294 7579 89602 7588
rect 86960 7404 87012 7410
rect 86960 7346 87012 7352
rect 86972 7206 87000 7346
rect 86960 7200 87012 7206
rect 86960 7142 87012 7148
rect 86972 6322 87000 7142
rect 89294 6556 89602 6565
rect 89294 6554 89300 6556
rect 89356 6554 89380 6556
rect 89436 6554 89460 6556
rect 89516 6554 89540 6556
rect 89596 6554 89602 6556
rect 89356 6502 89358 6554
rect 89538 6502 89540 6554
rect 89294 6500 89300 6502
rect 89356 6500 89380 6502
rect 89436 6500 89460 6502
rect 89516 6500 89540 6502
rect 89596 6500 89602 6502
rect 89294 6491 89602 6500
rect 86960 6316 87012 6322
rect 86960 6258 87012 6264
rect 87236 6112 87288 6118
rect 87236 6054 87288 6060
rect 87248 3058 87276 6054
rect 89294 5468 89602 5477
rect 89294 5466 89300 5468
rect 89356 5466 89380 5468
rect 89436 5466 89460 5468
rect 89516 5466 89540 5468
rect 89596 5466 89602 5468
rect 89356 5414 89358 5466
rect 89538 5414 89540 5466
rect 89294 5412 89300 5414
rect 89356 5412 89380 5414
rect 89436 5412 89460 5414
rect 89516 5412 89540 5414
rect 89596 5412 89602 5414
rect 89294 5403 89602 5412
rect 89294 4380 89602 4389
rect 89294 4378 89300 4380
rect 89356 4378 89380 4380
rect 89436 4378 89460 4380
rect 89516 4378 89540 4380
rect 89596 4378 89602 4380
rect 89356 4326 89358 4378
rect 89538 4326 89540 4378
rect 89294 4324 89300 4326
rect 89356 4324 89380 4326
rect 89436 4324 89460 4326
rect 89516 4324 89540 4326
rect 89596 4324 89602 4326
rect 89294 4315 89602 4324
rect 89294 3292 89602 3301
rect 89294 3290 89300 3292
rect 89356 3290 89380 3292
rect 89436 3290 89460 3292
rect 89516 3290 89540 3292
rect 89596 3290 89602 3292
rect 89356 3238 89358 3290
rect 89538 3238 89540 3290
rect 89294 3236 89300 3238
rect 89356 3236 89380 3238
rect 89436 3236 89460 3238
rect 89516 3236 89540 3238
rect 89596 3236 89602 3238
rect 89294 3227 89602 3236
rect 87236 3052 87288 3058
rect 87236 2994 87288 3000
rect 89168 2916 89220 2922
rect 89168 2858 89220 2864
rect 86960 2848 87012 2854
rect 86960 2790 87012 2796
rect 86500 1420 86552 1426
rect 86500 1362 86552 1368
rect 86592 1420 86644 1426
rect 86592 1362 86644 1368
rect 86512 1222 86540 1362
rect 86500 1216 86552 1222
rect 86500 1158 86552 1164
rect 86972 800 87000 2790
rect 89180 2446 89208 2858
rect 89534 2544 89590 2553
rect 89534 2479 89536 2488
rect 89588 2479 89590 2488
rect 89536 2450 89588 2456
rect 87604 2440 87656 2446
rect 87604 2382 87656 2388
rect 87696 2440 87748 2446
rect 87696 2382 87748 2388
rect 88984 2440 89036 2446
rect 88984 2382 89036 2388
rect 89168 2440 89220 2446
rect 89168 2382 89220 2388
rect 90456 2440 90508 2446
rect 90456 2382 90508 2388
rect 87616 800 87644 2382
rect 87708 1154 87736 2382
rect 88248 2304 88300 2310
rect 88248 2246 88300 2252
rect 87696 1148 87748 1154
rect 87696 1090 87748 1096
rect 88260 800 88288 2246
rect 88996 1465 89024 2382
rect 89168 2304 89220 2310
rect 89168 2246 89220 2252
rect 90180 2304 90232 2310
rect 90180 2246 90232 2252
rect 88982 1456 89038 1465
rect 88982 1391 89038 1400
rect 83844 734 84056 762
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 89180 762 89208 2246
rect 89294 2204 89602 2213
rect 89294 2202 89300 2204
rect 89356 2202 89380 2204
rect 89436 2202 89460 2204
rect 89516 2202 89540 2204
rect 89596 2202 89602 2204
rect 89356 2150 89358 2202
rect 89538 2150 89540 2202
rect 89294 2148 89300 2150
rect 89356 2148 89380 2150
rect 89436 2148 89460 2150
rect 89516 2148 89540 2150
rect 89596 2148 89602 2150
rect 89294 2139 89602 2148
rect 89718 2136 89774 2145
rect 89718 2071 89774 2080
rect 89442 1864 89498 1873
rect 89442 1799 89498 1808
rect 89536 1828 89588 1834
rect 89352 1488 89404 1494
rect 89350 1456 89352 1465
rect 89404 1456 89406 1465
rect 89456 1426 89484 1799
rect 89536 1770 89588 1776
rect 89628 1828 89680 1834
rect 89628 1770 89680 1776
rect 89548 1544 89576 1770
rect 89640 1737 89668 1770
rect 89626 1728 89682 1737
rect 89626 1663 89682 1672
rect 89732 1562 89760 2071
rect 89810 1864 89866 1873
rect 89810 1799 89866 1808
rect 89824 1562 89852 1799
rect 89628 1556 89680 1562
rect 89548 1516 89628 1544
rect 89628 1498 89680 1504
rect 89720 1556 89772 1562
rect 89720 1498 89772 1504
rect 89812 1556 89864 1562
rect 89812 1498 89864 1504
rect 89350 1391 89406 1400
rect 89444 1420 89496 1426
rect 89444 1362 89496 1368
rect 89536 1420 89588 1426
rect 89536 1362 89588 1368
rect 89548 1222 89576 1362
rect 89536 1216 89588 1222
rect 89536 1158 89588 1164
rect 89456 870 89576 898
rect 89456 762 89484 870
rect 89548 800 89576 870
rect 90192 800 90220 2246
rect 90468 1290 90496 2382
rect 90928 1465 90956 26726
rect 91020 23730 91048 27270
rect 91388 26994 91416 27474
rect 91480 27470 91508 29200
rect 91468 27464 91520 27470
rect 91468 27406 91520 27412
rect 91928 27328 91980 27334
rect 91928 27270 91980 27276
rect 92202 27296 92258 27305
rect 91376 26988 91428 26994
rect 91376 26930 91428 26936
rect 91744 26920 91796 26926
rect 91742 26888 91744 26897
rect 91796 26888 91798 26897
rect 91742 26823 91798 26832
rect 91836 26852 91888 26858
rect 91836 26794 91888 26800
rect 91744 26784 91796 26790
rect 91744 26726 91796 26732
rect 91756 26450 91784 26726
rect 91744 26444 91796 26450
rect 91744 26386 91796 26392
rect 91848 26314 91876 26794
rect 91836 26308 91888 26314
rect 91836 26250 91888 26256
rect 91008 23724 91060 23730
rect 91008 23666 91060 23672
rect 91940 10606 91968 27270
rect 92202 27231 92258 27240
rect 92216 26858 92244 27231
rect 92400 27112 92428 29294
rect 93398 29294 93532 29322
rect 93398 29200 93454 29294
rect 92756 27396 92808 27402
rect 92756 27338 92808 27344
rect 92480 27124 92532 27130
rect 92400 27084 92480 27112
rect 92480 27066 92532 27072
rect 92204 26852 92256 26858
rect 92204 26794 92256 26800
rect 92768 26625 92796 27338
rect 92848 27328 92900 27334
rect 92848 27270 92900 27276
rect 92754 26616 92810 26625
rect 92754 26551 92810 26560
rect 92860 26489 92888 27270
rect 92846 26480 92902 26489
rect 92846 26415 92902 26424
rect 93504 26246 93532 29294
rect 94042 29200 94098 30000
rect 94686 29322 94742 30000
rect 94686 29294 95188 29322
rect 94686 29200 94742 29294
rect 93676 27872 93728 27878
rect 93676 27814 93728 27820
rect 93688 26382 93716 27814
rect 94056 26858 94084 29200
rect 94872 27532 94924 27538
rect 94872 27474 94924 27480
rect 94596 27464 94648 27470
rect 94596 27406 94648 27412
rect 94884 27418 94912 27474
rect 94412 27328 94464 27334
rect 94412 27270 94464 27276
rect 94424 27062 94452 27270
rect 94608 27062 94636 27406
rect 94884 27390 95004 27418
rect 94688 27328 94740 27334
rect 94688 27270 94740 27276
rect 94872 27328 94924 27334
rect 94872 27270 94924 27276
rect 94412 27056 94464 27062
rect 94412 26998 94464 27004
rect 94596 27056 94648 27062
rect 94596 26998 94648 27004
rect 94044 26852 94096 26858
rect 94044 26794 94096 26800
rect 93676 26376 93728 26382
rect 93676 26318 93728 26324
rect 93492 26240 93544 26246
rect 93492 26182 93544 26188
rect 94700 25770 94728 27270
rect 94884 26994 94912 27270
rect 94872 26988 94924 26994
rect 94872 26930 94924 26936
rect 94688 25764 94740 25770
rect 94688 25706 94740 25712
rect 94780 22636 94832 22642
rect 94780 22578 94832 22584
rect 91928 10600 91980 10606
rect 91928 10542 91980 10548
rect 92202 2544 92258 2553
rect 92202 2479 92258 2488
rect 91468 2440 91520 2446
rect 91468 2382 91520 2388
rect 92112 2440 92164 2446
rect 92112 2382 92164 2388
rect 90914 1456 90970 1465
rect 90914 1391 90970 1400
rect 90456 1284 90508 1290
rect 90456 1226 90508 1232
rect 91480 800 91508 2382
rect 91560 2304 91612 2310
rect 91560 2246 91612 2252
rect 91572 1766 91600 2246
rect 91560 1760 91612 1766
rect 91560 1702 91612 1708
rect 92124 800 92152 2382
rect 92216 2310 92244 2479
rect 92756 2440 92808 2446
rect 92756 2382 92808 2388
rect 94320 2440 94372 2446
rect 94320 2382 94372 2388
rect 92296 2372 92348 2378
rect 92296 2314 92348 2320
rect 92204 2304 92256 2310
rect 92204 2246 92256 2252
rect 92308 2145 92336 2314
rect 92294 2136 92350 2145
rect 92294 2071 92350 2080
rect 92768 800 92796 2382
rect 93032 2304 93084 2310
rect 93032 2246 93084 2252
rect 94044 2304 94096 2310
rect 94044 2246 94096 2252
rect 93044 1358 93072 2246
rect 93032 1352 93084 1358
rect 93032 1294 93084 1300
rect 94056 800 94084 2246
rect 94332 1562 94360 2382
rect 94688 2372 94740 2378
rect 94688 2314 94740 2320
rect 94320 1556 94372 1562
rect 94320 1498 94372 1504
rect 94700 800 94728 2314
rect 94792 1834 94820 22578
rect 94976 22574 95004 27390
rect 95160 27112 95188 29294
rect 95974 29200 96030 30000
rect 96618 29322 96674 30000
rect 96618 29294 96936 29322
rect 96618 29200 96674 29294
rect 95988 27606 96016 29200
rect 96908 27606 96936 29294
rect 97906 29200 97962 30000
rect 98550 29200 98606 30000
rect 99838 29200 99894 30000
rect 100482 29322 100538 30000
rect 100482 29294 100616 29322
rect 100482 29200 100538 29294
rect 95792 27600 95844 27606
rect 95976 27600 96028 27606
rect 95792 27542 95844 27548
rect 95882 27568 95938 27577
rect 95804 27130 95832 27542
rect 96896 27600 96948 27606
rect 95976 27542 96028 27548
rect 96710 27568 96766 27577
rect 95882 27503 95938 27512
rect 96896 27542 96948 27548
rect 97920 27554 97948 29200
rect 98000 27600 98052 27606
rect 97920 27548 98000 27554
rect 97920 27542 98052 27548
rect 97920 27526 98040 27542
rect 98564 27538 98592 29200
rect 99852 27606 99880 29200
rect 99840 27600 99892 27606
rect 99840 27542 99892 27548
rect 98552 27532 98604 27538
rect 96710 27503 96766 27512
rect 95240 27124 95292 27130
rect 95160 27084 95240 27112
rect 95240 27066 95292 27072
rect 95792 27124 95844 27130
rect 95792 27066 95844 27072
rect 95896 26994 95924 27503
rect 96724 27470 96752 27503
rect 98552 27474 98604 27480
rect 96712 27464 96764 27470
rect 96250 27432 96306 27441
rect 96712 27406 96764 27412
rect 98184 27464 98236 27470
rect 98184 27406 98236 27412
rect 99380 27464 99432 27470
rect 99380 27406 99432 27412
rect 99564 27464 99616 27470
rect 99564 27406 99616 27412
rect 96250 27367 96306 27376
rect 96436 27396 96488 27402
rect 96264 27334 96292 27367
rect 96436 27338 96488 27344
rect 97172 27396 97224 27402
rect 97172 27338 97224 27344
rect 96252 27328 96304 27334
rect 96448 27305 96476 27338
rect 96712 27328 96764 27334
rect 96252 27270 96304 27276
rect 96434 27296 96490 27305
rect 96434 27231 96490 27240
rect 96710 27296 96712 27305
rect 96764 27296 96766 27305
rect 96710 27231 96766 27240
rect 97184 27169 97212 27338
rect 97170 27160 97226 27169
rect 97170 27095 97226 27104
rect 95240 26988 95292 26994
rect 95240 26930 95292 26936
rect 95884 26988 95936 26994
rect 95884 26930 95936 26936
rect 95976 26988 96028 26994
rect 95976 26930 96028 26936
rect 94964 22568 95016 22574
rect 94964 22510 95016 22516
rect 94976 14958 95004 22510
rect 94964 14952 95016 14958
rect 94964 14894 95016 14900
rect 95252 11898 95280 26930
rect 95790 26616 95846 26625
rect 95790 26551 95846 26560
rect 95804 26518 95832 26551
rect 95792 26512 95844 26518
rect 95792 26454 95844 26460
rect 95988 26353 96016 26930
rect 95974 26344 96030 26353
rect 95974 26279 96030 26288
rect 98196 22778 98224 27406
rect 98184 22772 98236 22778
rect 98184 22714 98236 22720
rect 99392 12646 99420 27406
rect 99576 27130 99604 27406
rect 100588 27130 100616 29294
rect 101126 29200 101182 30000
rect 102414 29322 102470 30000
rect 103058 29322 103114 30000
rect 104346 29322 104402 30000
rect 104990 29322 105046 30000
rect 102414 29294 102732 29322
rect 102414 29200 102470 29294
rect 100944 27600 100996 27606
rect 100944 27542 100996 27548
rect 100956 27402 100984 27542
rect 101140 27470 101168 29200
rect 101680 27668 101732 27674
rect 101680 27610 101732 27616
rect 101128 27464 101180 27470
rect 101128 27406 101180 27412
rect 100944 27396 100996 27402
rect 100944 27338 100996 27344
rect 99564 27124 99616 27130
rect 99564 27066 99616 27072
rect 100576 27124 100628 27130
rect 100576 27066 100628 27072
rect 101692 27062 101720 27610
rect 102704 27470 102732 29294
rect 103058 29294 103192 29322
rect 103058 29200 103114 29294
rect 103164 27606 103192 29294
rect 104346 29294 104664 29322
rect 104346 29200 104402 29294
rect 104018 27772 104326 27781
rect 104018 27770 104024 27772
rect 104080 27770 104104 27772
rect 104160 27770 104184 27772
rect 104240 27770 104264 27772
rect 104320 27770 104326 27772
rect 104080 27718 104082 27770
rect 104262 27718 104264 27770
rect 104018 27716 104024 27718
rect 104080 27716 104104 27718
rect 104160 27716 104184 27718
rect 104240 27716 104264 27718
rect 104320 27716 104326 27718
rect 104018 27707 104326 27716
rect 103152 27600 103204 27606
rect 103152 27542 103204 27548
rect 102692 27464 102744 27470
rect 102692 27406 102744 27412
rect 102784 27464 102836 27470
rect 102784 27406 102836 27412
rect 101680 27056 101732 27062
rect 101680 26998 101732 27004
rect 100852 26988 100904 26994
rect 100852 26930 100904 26936
rect 100206 26888 100262 26897
rect 100206 26823 100208 26832
rect 100260 26823 100262 26832
rect 100208 26794 100260 26800
rect 100864 26586 100892 26930
rect 100852 26580 100904 26586
rect 100852 26522 100904 26528
rect 102796 26450 102824 27406
rect 104636 27130 104664 29294
rect 104990 29294 105400 29322
rect 104990 29200 105046 29294
rect 105372 27470 105400 29294
rect 105634 29200 105690 30000
rect 106922 29200 106978 30000
rect 107566 29200 107622 30000
rect 108854 29322 108910 30000
rect 109498 29322 109554 30000
rect 110786 29322 110842 30000
rect 111430 29322 111486 30000
rect 108854 29294 108988 29322
rect 108854 29200 108910 29294
rect 105648 27606 105676 29200
rect 105636 27600 105688 27606
rect 105636 27542 105688 27548
rect 106936 27470 106964 29200
rect 107580 27588 107608 29200
rect 107660 27600 107712 27606
rect 107580 27560 107660 27588
rect 108960 27588 108988 29294
rect 109498 29294 109816 29322
rect 109498 29200 109554 29294
rect 109040 27600 109092 27606
rect 108960 27560 109040 27588
rect 107660 27542 107712 27548
rect 109040 27542 109092 27548
rect 109788 27470 109816 29294
rect 110786 29294 111104 29322
rect 110786 29200 110842 29294
rect 110972 27532 111024 27538
rect 110972 27474 111024 27480
rect 105360 27464 105412 27470
rect 104990 27432 105046 27441
rect 104716 27396 104768 27402
rect 105360 27406 105412 27412
rect 106372 27464 106424 27470
rect 106372 27406 106424 27412
rect 106924 27464 106976 27470
rect 106924 27406 106976 27412
rect 108488 27464 108540 27470
rect 108488 27406 108540 27412
rect 109592 27464 109644 27470
rect 109592 27406 109644 27412
rect 109776 27464 109828 27470
rect 109776 27406 109828 27412
rect 104990 27367 104992 27376
rect 104716 27338 104768 27344
rect 105044 27367 105046 27376
rect 104992 27338 105044 27344
rect 104624 27124 104676 27130
rect 104624 27066 104676 27072
rect 104728 27062 104756 27338
rect 104808 27328 104860 27334
rect 104808 27270 104860 27276
rect 104900 27328 104952 27334
rect 105636 27328 105688 27334
rect 104900 27270 104952 27276
rect 105634 27296 105636 27305
rect 105688 27296 105690 27305
rect 104716 27056 104768 27062
rect 104716 26998 104768 27004
rect 103336 26988 103388 26994
rect 103336 26930 103388 26936
rect 103348 26518 103376 26930
rect 104348 26920 104400 26926
rect 104820 26897 104848 27270
rect 104912 27033 104940 27270
rect 105634 27231 105690 27240
rect 104898 27024 104954 27033
rect 104898 26959 104954 26968
rect 105544 26988 105596 26994
rect 105544 26930 105596 26936
rect 104348 26862 104400 26868
rect 104806 26888 104862 26897
rect 104018 26684 104326 26693
rect 104018 26682 104024 26684
rect 104080 26682 104104 26684
rect 104160 26682 104184 26684
rect 104240 26682 104264 26684
rect 104320 26682 104326 26684
rect 104080 26630 104082 26682
rect 104262 26630 104264 26682
rect 104018 26628 104024 26630
rect 104080 26628 104104 26630
rect 104160 26628 104184 26630
rect 104240 26628 104264 26630
rect 104320 26628 104326 26630
rect 104018 26619 104326 26628
rect 104360 26586 104388 26862
rect 104806 26823 104862 26832
rect 104900 26852 104952 26858
rect 104900 26794 104952 26800
rect 104348 26580 104400 26586
rect 104348 26522 104400 26528
rect 103336 26512 103388 26518
rect 103336 26454 103388 26460
rect 102784 26444 102836 26450
rect 102784 26386 102836 26392
rect 102232 24132 102284 24138
rect 102232 24074 102284 24080
rect 99380 12640 99432 12646
rect 99380 12582 99432 12588
rect 95240 11892 95292 11898
rect 95240 11834 95292 11840
rect 99656 11824 99708 11830
rect 99656 11766 99708 11772
rect 97816 3596 97868 3602
rect 97816 3538 97868 3544
rect 96620 2372 96672 2378
rect 96620 2314 96672 2320
rect 94964 2304 95016 2310
rect 94964 2246 95016 2252
rect 95976 2304 96028 2310
rect 95976 2246 96028 2252
rect 94780 1828 94832 1834
rect 94780 1770 94832 1776
rect 94976 1494 95004 2246
rect 94964 1488 95016 1494
rect 94964 1430 95016 1436
rect 95988 800 96016 2246
rect 96632 800 96660 2314
rect 97080 2304 97132 2310
rect 97080 2246 97132 2252
rect 97092 1426 97120 2246
rect 97828 1562 97856 3538
rect 98552 2848 98604 2854
rect 98552 2790 98604 2796
rect 97908 2372 97960 2378
rect 97908 2314 97960 2320
rect 97816 1556 97868 1562
rect 97816 1498 97868 1504
rect 97080 1420 97132 1426
rect 97080 1362 97132 1368
rect 97920 800 97948 2314
rect 98184 2304 98236 2310
rect 98184 2246 98236 2252
rect 98196 1698 98224 2246
rect 98184 1692 98236 1698
rect 98184 1634 98236 1640
rect 98564 800 98592 2790
rect 99668 2446 99696 11766
rect 101496 3460 101548 3466
rect 101496 3402 101548 3408
rect 101508 3058 101536 3402
rect 101496 3052 101548 3058
rect 101496 2994 101548 3000
rect 102244 2650 102272 24074
rect 102692 19508 102744 19514
rect 102692 19450 102744 19456
rect 102704 3058 102732 19450
rect 102784 3188 102836 3194
rect 102784 3130 102836 3136
rect 102796 3058 102824 3130
rect 102692 3052 102744 3058
rect 102692 2994 102744 3000
rect 102784 3052 102836 3058
rect 102784 2994 102836 3000
rect 102416 2848 102468 2854
rect 102416 2790 102468 2796
rect 102232 2644 102284 2650
rect 102232 2586 102284 2592
rect 99656 2440 99708 2446
rect 99656 2382 99708 2388
rect 100484 2440 100536 2446
rect 100484 2382 100536 2388
rect 100668 2440 100720 2446
rect 100668 2382 100720 2388
rect 99196 2372 99248 2378
rect 99196 2314 99248 2320
rect 99208 800 99236 2314
rect 100496 800 100524 2382
rect 100680 1766 100708 2382
rect 101128 2372 101180 2378
rect 101128 2314 101180 2320
rect 100852 1828 100904 1834
rect 100852 1770 100904 1776
rect 100668 1760 100720 1766
rect 100668 1702 100720 1708
rect 100864 1562 100892 1770
rect 100852 1556 100904 1562
rect 100852 1498 100904 1504
rect 101140 800 101168 2314
rect 102428 800 102456 2790
rect 103348 2650 103376 26454
rect 104018 25596 104326 25605
rect 104018 25594 104024 25596
rect 104080 25594 104104 25596
rect 104160 25594 104184 25596
rect 104240 25594 104264 25596
rect 104320 25594 104326 25596
rect 104080 25542 104082 25594
rect 104262 25542 104264 25594
rect 104018 25540 104024 25542
rect 104080 25540 104104 25542
rect 104160 25540 104184 25542
rect 104240 25540 104264 25542
rect 104320 25540 104326 25542
rect 104018 25531 104326 25540
rect 104018 24508 104326 24517
rect 104018 24506 104024 24508
rect 104080 24506 104104 24508
rect 104160 24506 104184 24508
rect 104240 24506 104264 24508
rect 104320 24506 104326 24508
rect 104080 24454 104082 24506
rect 104262 24454 104264 24506
rect 104018 24452 104024 24454
rect 104080 24452 104104 24454
rect 104160 24452 104184 24454
rect 104240 24452 104264 24454
rect 104320 24452 104326 24454
rect 104018 24443 104326 24452
rect 104018 23420 104326 23429
rect 104018 23418 104024 23420
rect 104080 23418 104104 23420
rect 104160 23418 104184 23420
rect 104240 23418 104264 23420
rect 104320 23418 104326 23420
rect 104080 23366 104082 23418
rect 104262 23366 104264 23418
rect 104018 23364 104024 23366
rect 104080 23364 104104 23366
rect 104160 23364 104184 23366
rect 104240 23364 104264 23366
rect 104320 23364 104326 23366
rect 104018 23355 104326 23364
rect 104018 22332 104326 22341
rect 104018 22330 104024 22332
rect 104080 22330 104104 22332
rect 104160 22330 104184 22332
rect 104240 22330 104264 22332
rect 104320 22330 104326 22332
rect 104080 22278 104082 22330
rect 104262 22278 104264 22330
rect 104018 22276 104024 22278
rect 104080 22276 104104 22278
rect 104160 22276 104184 22278
rect 104240 22276 104264 22278
rect 104320 22276 104326 22278
rect 104018 22267 104326 22276
rect 104018 21244 104326 21253
rect 104018 21242 104024 21244
rect 104080 21242 104104 21244
rect 104160 21242 104184 21244
rect 104240 21242 104264 21244
rect 104320 21242 104326 21244
rect 104080 21190 104082 21242
rect 104262 21190 104264 21242
rect 104018 21188 104024 21190
rect 104080 21188 104104 21190
rect 104160 21188 104184 21190
rect 104240 21188 104264 21190
rect 104320 21188 104326 21190
rect 104018 21179 104326 21188
rect 104018 20156 104326 20165
rect 104018 20154 104024 20156
rect 104080 20154 104104 20156
rect 104160 20154 104184 20156
rect 104240 20154 104264 20156
rect 104320 20154 104326 20156
rect 104080 20102 104082 20154
rect 104262 20102 104264 20154
rect 104018 20100 104024 20102
rect 104080 20100 104104 20102
rect 104160 20100 104184 20102
rect 104240 20100 104264 20102
rect 104320 20100 104326 20102
rect 104018 20091 104326 20100
rect 104018 19068 104326 19077
rect 104018 19066 104024 19068
rect 104080 19066 104104 19068
rect 104160 19066 104184 19068
rect 104240 19066 104264 19068
rect 104320 19066 104326 19068
rect 104080 19014 104082 19066
rect 104262 19014 104264 19066
rect 104018 19012 104024 19014
rect 104080 19012 104104 19014
rect 104160 19012 104184 19014
rect 104240 19012 104264 19014
rect 104320 19012 104326 19014
rect 104018 19003 104326 19012
rect 104018 17980 104326 17989
rect 104018 17978 104024 17980
rect 104080 17978 104104 17980
rect 104160 17978 104184 17980
rect 104240 17978 104264 17980
rect 104320 17978 104326 17980
rect 104080 17926 104082 17978
rect 104262 17926 104264 17978
rect 104018 17924 104024 17926
rect 104080 17924 104104 17926
rect 104160 17924 104184 17926
rect 104240 17924 104264 17926
rect 104320 17924 104326 17926
rect 104018 17915 104326 17924
rect 104018 16892 104326 16901
rect 104018 16890 104024 16892
rect 104080 16890 104104 16892
rect 104160 16890 104184 16892
rect 104240 16890 104264 16892
rect 104320 16890 104326 16892
rect 104080 16838 104082 16890
rect 104262 16838 104264 16890
rect 104018 16836 104024 16838
rect 104080 16836 104104 16838
rect 104160 16836 104184 16838
rect 104240 16836 104264 16838
rect 104320 16836 104326 16838
rect 104018 16827 104326 16836
rect 104018 15804 104326 15813
rect 104018 15802 104024 15804
rect 104080 15802 104104 15804
rect 104160 15802 104184 15804
rect 104240 15802 104264 15804
rect 104320 15802 104326 15804
rect 104080 15750 104082 15802
rect 104262 15750 104264 15802
rect 104018 15748 104024 15750
rect 104080 15748 104104 15750
rect 104160 15748 104184 15750
rect 104240 15748 104264 15750
rect 104320 15748 104326 15750
rect 104018 15739 104326 15748
rect 104018 14716 104326 14725
rect 104018 14714 104024 14716
rect 104080 14714 104104 14716
rect 104160 14714 104184 14716
rect 104240 14714 104264 14716
rect 104320 14714 104326 14716
rect 104080 14662 104082 14714
rect 104262 14662 104264 14714
rect 104018 14660 104024 14662
rect 104080 14660 104104 14662
rect 104160 14660 104184 14662
rect 104240 14660 104264 14662
rect 104320 14660 104326 14662
rect 104018 14651 104326 14660
rect 104018 13628 104326 13637
rect 104018 13626 104024 13628
rect 104080 13626 104104 13628
rect 104160 13626 104184 13628
rect 104240 13626 104264 13628
rect 104320 13626 104326 13628
rect 104080 13574 104082 13626
rect 104262 13574 104264 13626
rect 104018 13572 104024 13574
rect 104080 13572 104104 13574
rect 104160 13572 104184 13574
rect 104240 13572 104264 13574
rect 104320 13572 104326 13574
rect 104018 13563 104326 13572
rect 104018 12540 104326 12549
rect 104018 12538 104024 12540
rect 104080 12538 104104 12540
rect 104160 12538 104184 12540
rect 104240 12538 104264 12540
rect 104320 12538 104326 12540
rect 104080 12486 104082 12538
rect 104262 12486 104264 12538
rect 104018 12484 104024 12486
rect 104080 12484 104104 12486
rect 104160 12484 104184 12486
rect 104240 12484 104264 12486
rect 104320 12484 104326 12486
rect 104018 12475 104326 12484
rect 104018 11452 104326 11461
rect 104018 11450 104024 11452
rect 104080 11450 104104 11452
rect 104160 11450 104184 11452
rect 104240 11450 104264 11452
rect 104320 11450 104326 11452
rect 104080 11398 104082 11450
rect 104262 11398 104264 11450
rect 104018 11396 104024 11398
rect 104080 11396 104104 11398
rect 104160 11396 104184 11398
rect 104240 11396 104264 11398
rect 104320 11396 104326 11398
rect 104018 11387 104326 11396
rect 104018 10364 104326 10373
rect 104018 10362 104024 10364
rect 104080 10362 104104 10364
rect 104160 10362 104184 10364
rect 104240 10362 104264 10364
rect 104320 10362 104326 10364
rect 104080 10310 104082 10362
rect 104262 10310 104264 10362
rect 104018 10308 104024 10310
rect 104080 10308 104104 10310
rect 104160 10308 104184 10310
rect 104240 10308 104264 10310
rect 104320 10308 104326 10310
rect 104018 10299 104326 10308
rect 104018 9276 104326 9285
rect 104018 9274 104024 9276
rect 104080 9274 104104 9276
rect 104160 9274 104184 9276
rect 104240 9274 104264 9276
rect 104320 9274 104326 9276
rect 104080 9222 104082 9274
rect 104262 9222 104264 9274
rect 104018 9220 104024 9222
rect 104080 9220 104104 9222
rect 104160 9220 104184 9222
rect 104240 9220 104264 9222
rect 104320 9220 104326 9222
rect 104018 9211 104326 9220
rect 104018 8188 104326 8197
rect 104018 8186 104024 8188
rect 104080 8186 104104 8188
rect 104160 8186 104184 8188
rect 104240 8186 104264 8188
rect 104320 8186 104326 8188
rect 104080 8134 104082 8186
rect 104262 8134 104264 8186
rect 104018 8132 104024 8134
rect 104080 8132 104104 8134
rect 104160 8132 104184 8134
rect 104240 8132 104264 8134
rect 104320 8132 104326 8134
rect 104018 8123 104326 8132
rect 104018 7100 104326 7109
rect 104018 7098 104024 7100
rect 104080 7098 104104 7100
rect 104160 7098 104184 7100
rect 104240 7098 104264 7100
rect 104320 7098 104326 7100
rect 104080 7046 104082 7098
rect 104262 7046 104264 7098
rect 104018 7044 104024 7046
rect 104080 7044 104104 7046
rect 104160 7044 104184 7046
rect 104240 7044 104264 7046
rect 104320 7044 104326 7046
rect 104018 7035 104326 7044
rect 104018 6012 104326 6021
rect 104018 6010 104024 6012
rect 104080 6010 104104 6012
rect 104160 6010 104184 6012
rect 104240 6010 104264 6012
rect 104320 6010 104326 6012
rect 104080 5958 104082 6010
rect 104262 5958 104264 6010
rect 104018 5956 104024 5958
rect 104080 5956 104104 5958
rect 104160 5956 104184 5958
rect 104240 5956 104264 5958
rect 104320 5956 104326 5958
rect 104018 5947 104326 5956
rect 104018 4924 104326 4933
rect 104018 4922 104024 4924
rect 104080 4922 104104 4924
rect 104160 4922 104184 4924
rect 104240 4922 104264 4924
rect 104320 4922 104326 4924
rect 104080 4870 104082 4922
rect 104262 4870 104264 4922
rect 104018 4868 104024 4870
rect 104080 4868 104104 4870
rect 104160 4868 104184 4870
rect 104240 4868 104264 4870
rect 104320 4868 104326 4870
rect 104018 4859 104326 4868
rect 104018 3836 104326 3845
rect 104018 3834 104024 3836
rect 104080 3834 104104 3836
rect 104160 3834 104184 3836
rect 104240 3834 104264 3836
rect 104320 3834 104326 3836
rect 104080 3782 104082 3834
rect 104262 3782 104264 3834
rect 104018 3780 104024 3782
rect 104080 3780 104104 3782
rect 104160 3780 104184 3782
rect 104240 3780 104264 3782
rect 104320 3780 104326 3782
rect 104018 3771 104326 3780
rect 103992 3194 104296 3210
rect 103992 3188 104308 3194
rect 103992 3182 104256 3188
rect 103992 3126 104020 3182
rect 104256 3130 104308 3136
rect 103980 3120 104032 3126
rect 103980 3062 104032 3068
rect 104018 2748 104326 2757
rect 104018 2746 104024 2748
rect 104080 2746 104104 2748
rect 104160 2746 104184 2748
rect 104240 2746 104264 2748
rect 104320 2746 104326 2748
rect 104080 2694 104082 2746
rect 104262 2694 104264 2746
rect 104018 2692 104024 2694
rect 104080 2692 104104 2694
rect 104160 2692 104184 2694
rect 104240 2692 104264 2694
rect 104320 2692 104326 2694
rect 104018 2683 104326 2692
rect 103336 2644 103388 2650
rect 103336 2586 103388 2592
rect 104532 2644 104584 2650
rect 104532 2586 104584 2592
rect 104544 2446 104572 2586
rect 104912 2446 104940 26794
rect 105556 10538 105584 26930
rect 106384 21894 106412 27406
rect 108500 26926 108528 27406
rect 109604 26926 109632 27406
rect 110052 27328 110104 27334
rect 110052 27270 110104 27276
rect 110064 27130 110092 27270
rect 110052 27124 110104 27130
rect 110052 27066 110104 27072
rect 108488 26920 108540 26926
rect 108488 26862 108540 26868
rect 109592 26920 109644 26926
rect 109592 26862 109644 26868
rect 110984 26586 111012 27474
rect 111076 27470 111104 29294
rect 111430 29294 111564 29322
rect 111430 29200 111486 29294
rect 111064 27464 111116 27470
rect 111064 27406 111116 27412
rect 111536 27130 111564 29294
rect 112074 29200 112130 30000
rect 113362 29322 113418 30000
rect 114006 29322 114062 30000
rect 115294 29322 115350 30000
rect 115938 29322 115994 30000
rect 113362 29294 113680 29322
rect 113362 29200 113418 29294
rect 112088 27470 112116 29200
rect 113652 27606 113680 29294
rect 114006 29294 114508 29322
rect 114006 29200 114062 29294
rect 113640 27600 113692 27606
rect 113640 27542 113692 27548
rect 114480 27554 114508 29294
rect 115294 29294 115612 29322
rect 115294 29200 115350 29294
rect 115584 27606 115612 29294
rect 115938 29294 116072 29322
rect 115938 29200 115994 29294
rect 115572 27600 115624 27606
rect 114480 27526 114600 27554
rect 115572 27542 115624 27548
rect 114572 27470 114600 27526
rect 116044 27470 116072 29294
rect 117134 29200 117190 29209
rect 117226 29200 117282 30000
rect 117870 29200 117926 30000
rect 118514 29200 118570 30000
rect 119802 29200 119858 30000
rect 117134 29135 117190 29144
rect 117042 27976 117098 27985
rect 117042 27911 117098 27920
rect 116768 27532 116820 27538
rect 116768 27474 116820 27480
rect 112076 27464 112128 27470
rect 112076 27406 112128 27412
rect 114560 27464 114612 27470
rect 114560 27406 114612 27412
rect 116032 27464 116084 27470
rect 116032 27406 116084 27412
rect 112536 27328 112588 27334
rect 112536 27270 112588 27276
rect 114744 27328 114796 27334
rect 114744 27270 114796 27276
rect 115204 27328 115256 27334
rect 115204 27270 115256 27276
rect 111524 27124 111576 27130
rect 111524 27066 111576 27072
rect 111708 26988 111760 26994
rect 111708 26930 111760 26936
rect 110972 26580 111024 26586
rect 110972 26522 111024 26528
rect 107660 25288 107712 25294
rect 107660 25230 107712 25236
rect 106372 21888 106424 21894
rect 106372 21830 106424 21836
rect 105544 10532 105596 10538
rect 105544 10474 105596 10480
rect 107476 4140 107528 4146
rect 107476 4082 107528 4088
rect 107488 3126 107516 4082
rect 107476 3120 107528 3126
rect 107476 3062 107528 3068
rect 107488 2446 107516 3062
rect 107672 2922 107700 25230
rect 108120 13932 108172 13938
rect 108120 13874 108172 13880
rect 108132 12850 108160 13874
rect 108120 12844 108172 12850
rect 108120 12786 108172 12792
rect 107660 2916 107712 2922
rect 107660 2858 107712 2864
rect 108132 2446 108160 12786
rect 111720 10470 111748 26930
rect 112548 15366 112576 27270
rect 113640 26920 113692 26926
rect 113640 26862 113692 26868
rect 112536 15360 112588 15366
rect 112536 15302 112588 15308
rect 111708 10464 111760 10470
rect 111708 10406 111760 10412
rect 113652 10266 113680 26862
rect 114756 20466 114784 27270
rect 114744 20460 114796 20466
rect 114744 20402 114796 20408
rect 114756 19786 114784 20402
rect 114744 19780 114796 19786
rect 114744 19722 114796 19728
rect 113732 19712 113784 19718
rect 113732 19654 113784 19660
rect 113744 19514 113772 19654
rect 113732 19508 113784 19514
rect 113732 19450 113784 19456
rect 115216 17270 115244 27270
rect 116780 27062 116808 27474
rect 116768 27056 116820 27062
rect 116768 26998 116820 27004
rect 117056 26382 117084 27911
rect 117148 26994 117176 29135
rect 117240 27130 117268 29200
rect 117320 27464 117372 27470
rect 117320 27406 117372 27412
rect 117332 27305 117360 27406
rect 117318 27296 117374 27305
rect 117318 27231 117374 27240
rect 117228 27124 117280 27130
rect 117228 27066 117280 27072
rect 117136 26988 117188 26994
rect 117136 26930 117188 26936
rect 117780 26784 117832 26790
rect 117780 26726 117832 26732
rect 117412 26512 117464 26518
rect 117412 26454 117464 26460
rect 116860 26376 116912 26382
rect 116860 26318 116912 26324
rect 117044 26376 117096 26382
rect 117044 26318 117096 26324
rect 115940 20936 115992 20942
rect 115940 20878 115992 20884
rect 115952 20602 115980 20878
rect 115940 20596 115992 20602
rect 115940 20538 115992 20544
rect 115204 17264 115256 17270
rect 115204 17206 115256 17212
rect 113640 10260 113692 10266
rect 113640 10202 113692 10208
rect 115940 10056 115992 10062
rect 115940 9998 115992 10004
rect 114744 9988 114796 9994
rect 114744 9930 114796 9936
rect 114756 9586 114784 9930
rect 115388 9648 115440 9654
rect 115388 9590 115440 9596
rect 114744 9580 114796 9586
rect 114744 9522 114796 9528
rect 113640 8968 113692 8974
rect 113640 8910 113692 8916
rect 110052 6180 110104 6186
rect 110052 6122 110104 6128
rect 109776 3120 109828 3126
rect 109776 3062 109828 3068
rect 109500 2916 109552 2922
rect 109500 2858 109552 2864
rect 104532 2440 104584 2446
rect 104532 2382 104584 2388
rect 104900 2440 104952 2446
rect 104900 2382 104952 2388
rect 106004 2440 106056 2446
rect 106004 2382 106056 2388
rect 107476 2440 107528 2446
rect 107476 2382 107528 2388
rect 108120 2440 108172 2446
rect 108120 2382 108172 2388
rect 108304 2440 108356 2446
rect 108304 2382 108356 2388
rect 103060 2372 103112 2378
rect 103060 2314 103112 2320
rect 104992 2372 105044 2378
rect 104992 2314 105044 2320
rect 103072 800 103100 2314
rect 104348 2304 104400 2310
rect 104348 2246 104400 2252
rect 104360 800 104388 2246
rect 105004 800 105032 2314
rect 105268 2304 105320 2310
rect 105268 2246 105320 2252
rect 105636 2304 105688 2310
rect 105636 2246 105688 2252
rect 105280 1970 105308 2246
rect 105268 1964 105320 1970
rect 105268 1906 105320 1912
rect 105648 800 105676 2246
rect 106016 1834 106044 2382
rect 106924 2304 106976 2310
rect 106924 2246 106976 2252
rect 106004 1828 106056 1834
rect 106004 1770 106056 1776
rect 106936 800 106964 2246
rect 108316 1426 108344 2382
rect 108856 2372 108908 2378
rect 108856 2314 108908 2320
rect 107568 1420 107620 1426
rect 107568 1362 107620 1368
rect 108304 1420 108356 1426
rect 108304 1362 108356 1368
rect 107580 800 107608 1362
rect 108868 800 108896 2314
rect 109512 800 109540 2858
rect 109788 2854 109816 3062
rect 109776 2848 109828 2854
rect 109776 2790 109828 2796
rect 109788 1902 109816 2790
rect 110064 2514 110092 6122
rect 110236 3052 110288 3058
rect 110236 2994 110288 3000
rect 111432 3052 111484 3058
rect 111432 2994 111484 3000
rect 110248 2922 110276 2994
rect 110236 2916 110288 2922
rect 110236 2858 110288 2864
rect 110052 2508 110104 2514
rect 110052 2450 110104 2456
rect 110788 2440 110840 2446
rect 110788 2382 110840 2388
rect 109960 2304 110012 2310
rect 109960 2246 110012 2252
rect 109776 1896 109828 1902
rect 109776 1838 109828 1844
rect 109972 1630 110000 2246
rect 109960 1624 110012 1630
rect 109960 1566 110012 1572
rect 110800 800 110828 2382
rect 111444 800 111472 2994
rect 113652 2446 113680 8910
rect 114756 2650 114784 9522
rect 115400 8945 115428 9590
rect 115952 9450 115980 9998
rect 115940 9444 115992 9450
rect 115940 9386 115992 9392
rect 115386 8936 115442 8945
rect 115386 8871 115442 8880
rect 116216 7812 116268 7818
rect 116216 7754 116268 7760
rect 115664 5228 115716 5234
rect 115664 5170 115716 5176
rect 115676 4554 115704 5170
rect 115664 4548 115716 4554
rect 115664 4490 115716 4496
rect 116228 3058 116256 7754
rect 116872 4146 116900 26318
rect 117228 23656 117280 23662
rect 117228 23598 117280 23604
rect 117240 23225 117268 23598
rect 117226 23216 117282 23225
rect 117226 23151 117282 23160
rect 117320 21480 117372 21486
rect 117320 21422 117372 21428
rect 117332 21185 117360 21422
rect 117318 21176 117374 21185
rect 117318 21111 117374 21120
rect 117228 16584 117280 16590
rect 117228 16526 117280 16532
rect 117240 16425 117268 16526
rect 117226 16416 117282 16425
rect 117226 16351 117282 16360
rect 117424 15434 117452 26454
rect 117792 26314 117820 26726
rect 117780 26308 117832 26314
rect 117780 26250 117832 26256
rect 117884 25906 117912 29200
rect 117964 26988 118016 26994
rect 117964 26930 118016 26936
rect 117976 26625 118004 26930
rect 117962 26616 118018 26625
rect 117962 26551 118018 26560
rect 118528 26382 118556 29200
rect 118516 26376 118568 26382
rect 118516 26318 118568 26324
rect 118056 26308 118108 26314
rect 118056 26250 118108 26256
rect 117872 25900 117924 25906
rect 117872 25842 117924 25848
rect 117962 25256 118018 25265
rect 117962 25191 118018 25200
rect 117976 25158 118004 25191
rect 117964 25152 118016 25158
rect 117964 25094 118016 25100
rect 117964 24608 118016 24614
rect 117962 24576 117964 24585
rect 118016 24576 118018 24585
rect 117962 24511 118018 24520
rect 117962 22536 118018 22545
rect 117962 22471 117964 22480
rect 118016 22471 118018 22480
rect 117964 22442 118016 22448
rect 117596 21480 117648 21486
rect 117596 21422 117648 21428
rect 117608 21078 117636 21422
rect 117596 21072 117648 21078
rect 117596 21014 117648 21020
rect 118068 20874 118096 26250
rect 119816 25974 119844 29200
rect 119804 25968 119856 25974
rect 119804 25910 119856 25916
rect 118056 20868 118108 20874
rect 118056 20810 118108 20816
rect 117964 20800 118016 20806
rect 117964 20742 118016 20748
rect 117976 20505 118004 20742
rect 117962 20496 118018 20505
rect 117962 20431 118018 20440
rect 117962 19816 118018 19825
rect 117962 19751 118018 19760
rect 117976 19718 118004 19751
rect 117964 19712 118016 19718
rect 117964 19654 118016 19660
rect 117872 18760 117924 18766
rect 117872 18702 117924 18708
rect 117884 18465 117912 18702
rect 117964 18624 118016 18630
rect 117964 18566 118016 18572
rect 117870 18456 117926 18465
rect 117870 18391 117926 18400
rect 117872 18284 117924 18290
rect 117872 18226 117924 18232
rect 117688 18080 117740 18086
rect 117688 18022 117740 18028
rect 117412 15428 117464 15434
rect 117412 15370 117464 15376
rect 117320 11688 117372 11694
rect 117318 11656 117320 11665
rect 117412 11688 117464 11694
rect 117372 11656 117374 11665
rect 117412 11630 117464 11636
rect 117318 11591 117374 11600
rect 116860 4140 116912 4146
rect 116860 4082 116912 4088
rect 117136 3732 117188 3738
rect 117136 3674 117188 3680
rect 116676 3392 116728 3398
rect 116676 3334 116728 3340
rect 116216 3052 116268 3058
rect 116216 2994 116268 3000
rect 115940 2848 115992 2854
rect 115940 2790 115992 2796
rect 114744 2644 114796 2650
rect 114744 2586 114796 2592
rect 112076 2440 112128 2446
rect 112076 2382 112128 2388
rect 112444 2440 112496 2446
rect 112444 2382 112496 2388
rect 113640 2440 113692 2446
rect 113640 2382 113692 2388
rect 114008 2440 114060 2446
rect 114008 2382 114060 2388
rect 115296 2440 115348 2446
rect 115296 2382 115348 2388
rect 115570 2408 115626 2417
rect 112088 800 112116 2382
rect 112456 1766 112484 2382
rect 113364 2304 113416 2310
rect 113364 2246 113416 2252
rect 112444 1760 112496 1766
rect 112444 1702 112496 1708
rect 113376 800 113404 2246
rect 114020 800 114048 2382
rect 115308 800 115336 2382
rect 115570 2343 115626 2352
rect 115584 2310 115612 2343
rect 115572 2304 115624 2310
rect 115572 2246 115624 2252
rect 115952 800 115980 2790
rect 116400 2372 116452 2378
rect 116400 2314 116452 2320
rect 116584 2372 116636 2378
rect 116584 2314 116636 2320
rect 116412 2145 116440 2314
rect 116492 2304 116544 2310
rect 116492 2246 116544 2252
rect 116398 2136 116454 2145
rect 116398 2071 116454 2080
rect 116504 2038 116532 2246
rect 116492 2032 116544 2038
rect 116492 1974 116544 1980
rect 116596 800 116624 2314
rect 116688 1465 116716 3334
rect 117148 3194 117176 3674
rect 117424 3534 117452 11630
rect 117700 3738 117728 18022
rect 117884 17785 117912 18226
rect 117870 17776 117926 17785
rect 117870 17711 117926 17720
rect 117872 14408 117924 14414
rect 117870 14376 117872 14385
rect 117924 14376 117926 14385
rect 117870 14311 117926 14320
rect 117872 13932 117924 13938
rect 117872 13874 117924 13880
rect 117884 13705 117912 13874
rect 117870 13696 117926 13705
rect 117870 13631 117926 13640
rect 117976 13274 118004 18566
rect 118148 15904 118200 15910
rect 118148 15846 118200 15852
rect 118160 15745 118188 15846
rect 118146 15736 118202 15745
rect 118146 15671 118202 15680
rect 118056 15156 118108 15162
rect 118056 15098 118108 15104
rect 118068 14618 118096 15098
rect 118056 14612 118108 14618
rect 118056 14554 118108 14560
rect 118240 14068 118292 14074
rect 118240 14010 118292 14016
rect 118148 13320 118200 13326
rect 117976 13246 118096 13274
rect 118148 13262 118200 13268
rect 117964 13184 118016 13190
rect 117964 13126 118016 13132
rect 117976 13025 118004 13126
rect 117962 13016 118018 13025
rect 117962 12951 118018 12960
rect 117964 11280 118016 11286
rect 117964 11222 118016 11228
rect 117976 10985 118004 11222
rect 117962 10976 118018 10985
rect 117962 10911 118018 10920
rect 117964 9920 118016 9926
rect 117964 9862 118016 9868
rect 117976 9625 118004 9862
rect 117962 9616 118018 9625
rect 117962 9551 118018 9560
rect 117964 8356 118016 8362
rect 117964 8298 118016 8304
rect 117976 8265 118004 8298
rect 117962 8256 118018 8265
rect 117962 8191 118018 8200
rect 117964 7404 118016 7410
rect 117964 7346 118016 7352
rect 117976 6905 118004 7346
rect 118068 6914 118096 13246
rect 118160 12646 118188 13262
rect 118148 12640 118200 12646
rect 118148 12582 118200 12588
rect 118148 11552 118200 11558
rect 118148 11494 118200 11500
rect 118160 11150 118188 11494
rect 118148 11144 118200 11150
rect 118148 11086 118200 11092
rect 117962 6896 118018 6905
rect 118068 6886 118188 6914
rect 117962 6831 118018 6840
rect 117872 6316 117924 6322
rect 117872 6258 117924 6264
rect 117884 6225 117912 6258
rect 117870 6216 117926 6225
rect 117870 6151 117926 6160
rect 117964 5024 118016 5030
rect 117964 4966 118016 4972
rect 117976 4865 118004 4966
rect 117962 4856 118018 4865
rect 117962 4791 118018 4800
rect 117780 4548 117832 4554
rect 117780 4490 117832 4496
rect 117792 4185 117820 4490
rect 117778 4176 117834 4185
rect 117778 4111 117834 4120
rect 117964 3936 118016 3942
rect 117964 3878 118016 3884
rect 118056 3936 118108 3942
rect 118056 3878 118108 3884
rect 117688 3732 117740 3738
rect 117688 3674 117740 3680
rect 117412 3528 117464 3534
rect 117412 3470 117464 3476
rect 117872 3528 117924 3534
rect 117872 3470 117924 3476
rect 117136 3188 117188 3194
rect 117136 3130 117188 3136
rect 117424 3058 117452 3470
rect 117412 3052 117464 3058
rect 117412 2994 117464 3000
rect 117780 3052 117832 3058
rect 117780 2994 117832 3000
rect 116674 1456 116730 1465
rect 116674 1391 116730 1400
rect 89180 734 89484 762
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92754 0 92810 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 100482 0 100538 800
rect 101126 0 101182 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 104346 0 104402 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106922 0 106978 800
rect 107566 0 107622 800
rect 108854 0 108910 800
rect 109498 0 109554 800
rect 110786 0 110842 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 115294 0 115350 800
rect 115938 0 115994 800
rect 116582 0 116638 800
rect 117792 105 117820 2994
rect 117884 2825 117912 3470
rect 117870 2816 117926 2825
rect 117870 2751 117926 2760
rect 117976 1986 118004 3878
rect 118068 2106 118096 3878
rect 118160 2446 118188 6886
rect 118252 2582 118280 14010
rect 119804 4208 119856 4214
rect 119804 4150 119856 4156
rect 118516 3120 118568 3126
rect 118516 3062 118568 3068
rect 118240 2576 118292 2582
rect 118240 2518 118292 2524
rect 118148 2440 118200 2446
rect 118148 2382 118200 2388
rect 118056 2100 118108 2106
rect 118056 2042 118108 2048
rect 117884 1958 118004 1986
rect 117884 800 117912 1958
rect 118528 800 118556 3062
rect 119816 800 119844 4150
rect 117778 96 117834 105
rect 117778 31 117834 40
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119802 0 119858 800
<< via2 >>
rect 1214 28600 1270 28656
rect 2778 27920 2834 27976
rect 1398 26560 1454 26616
rect 1398 25880 1454 25936
rect 1398 24520 1454 24576
rect 1398 23840 1454 23896
rect 1398 23160 1454 23216
rect 1398 21836 1400 21856
rect 1400 21836 1452 21856
rect 1452 21836 1454 21856
rect 1398 21800 1454 21836
rect 1398 21120 1454 21176
rect 1398 19760 1454 19816
rect 1398 18400 1454 18456
rect 1398 17060 1454 17096
rect 1398 17040 1400 17060
rect 1400 17040 1452 17060
rect 1452 17040 1454 17060
rect 1398 15000 1454 15056
rect 1398 14320 1454 14376
rect 1398 12280 1454 12336
rect 1582 16360 1638 16416
rect 1398 11620 1454 11656
rect 1398 11600 1400 11620
rect 1400 11600 1452 11620
rect 1452 11600 1454 11620
rect 1398 10240 1454 10296
rect 1398 8200 1454 8256
rect 1398 7520 1454 7576
rect 1398 6180 1454 6216
rect 1398 6160 1400 6180
rect 1400 6160 1452 6180
rect 1452 6160 1454 6180
rect 1398 4800 1454 4856
rect 1858 19080 1914 19136
rect 1858 12960 1914 13016
rect 1858 9560 1914 9616
rect 1858 5480 1914 5536
rect 1582 3476 1584 3496
rect 1584 3476 1636 3496
rect 1636 3476 1638 3496
rect 1582 3440 1638 3476
rect 1398 2760 1454 2816
rect 2778 1400 2834 1456
rect 14462 27240 14518 27296
rect 15680 27770 15736 27772
rect 15760 27770 15816 27772
rect 15840 27770 15896 27772
rect 15920 27770 15976 27772
rect 15680 27718 15726 27770
rect 15726 27718 15736 27770
rect 15760 27718 15790 27770
rect 15790 27718 15802 27770
rect 15802 27718 15816 27770
rect 15840 27718 15854 27770
rect 15854 27718 15866 27770
rect 15866 27718 15896 27770
rect 15920 27718 15930 27770
rect 15930 27718 15976 27770
rect 15680 27716 15736 27718
rect 15760 27716 15816 27718
rect 15840 27716 15896 27718
rect 15920 27716 15976 27718
rect 15198 26968 15254 27024
rect 16210 27240 16266 27296
rect 15680 26682 15736 26684
rect 15760 26682 15816 26684
rect 15840 26682 15896 26684
rect 15920 26682 15976 26684
rect 15680 26630 15726 26682
rect 15726 26630 15736 26682
rect 15760 26630 15790 26682
rect 15790 26630 15802 26682
rect 15802 26630 15816 26682
rect 15840 26630 15854 26682
rect 15854 26630 15866 26682
rect 15866 26630 15896 26682
rect 15920 26630 15930 26682
rect 15930 26630 15976 26682
rect 15680 26628 15736 26630
rect 15760 26628 15816 26630
rect 15840 26628 15896 26630
rect 15920 26628 15976 26630
rect 15680 25594 15736 25596
rect 15760 25594 15816 25596
rect 15840 25594 15896 25596
rect 15920 25594 15976 25596
rect 15680 25542 15726 25594
rect 15726 25542 15736 25594
rect 15760 25542 15790 25594
rect 15790 25542 15802 25594
rect 15802 25542 15816 25594
rect 15840 25542 15854 25594
rect 15854 25542 15866 25594
rect 15866 25542 15896 25594
rect 15920 25542 15930 25594
rect 15930 25542 15976 25594
rect 15680 25540 15736 25542
rect 15760 25540 15816 25542
rect 15840 25540 15896 25542
rect 15920 25540 15976 25542
rect 15680 24506 15736 24508
rect 15760 24506 15816 24508
rect 15840 24506 15896 24508
rect 15920 24506 15976 24508
rect 15680 24454 15726 24506
rect 15726 24454 15736 24506
rect 15760 24454 15790 24506
rect 15790 24454 15802 24506
rect 15802 24454 15816 24506
rect 15840 24454 15854 24506
rect 15854 24454 15866 24506
rect 15866 24454 15896 24506
rect 15920 24454 15930 24506
rect 15930 24454 15976 24506
rect 15680 24452 15736 24454
rect 15760 24452 15816 24454
rect 15840 24452 15896 24454
rect 15920 24452 15976 24454
rect 15680 23418 15736 23420
rect 15760 23418 15816 23420
rect 15840 23418 15896 23420
rect 15920 23418 15976 23420
rect 15680 23366 15726 23418
rect 15726 23366 15736 23418
rect 15760 23366 15790 23418
rect 15790 23366 15802 23418
rect 15802 23366 15816 23418
rect 15840 23366 15854 23418
rect 15854 23366 15866 23418
rect 15866 23366 15896 23418
rect 15920 23366 15930 23418
rect 15930 23366 15976 23418
rect 15680 23364 15736 23366
rect 15760 23364 15816 23366
rect 15840 23364 15896 23366
rect 15920 23364 15976 23366
rect 15680 22330 15736 22332
rect 15760 22330 15816 22332
rect 15840 22330 15896 22332
rect 15920 22330 15976 22332
rect 15680 22278 15726 22330
rect 15726 22278 15736 22330
rect 15760 22278 15790 22330
rect 15790 22278 15802 22330
rect 15802 22278 15816 22330
rect 15840 22278 15854 22330
rect 15854 22278 15866 22330
rect 15866 22278 15896 22330
rect 15920 22278 15930 22330
rect 15930 22278 15976 22330
rect 15680 22276 15736 22278
rect 15760 22276 15816 22278
rect 15840 22276 15896 22278
rect 15920 22276 15976 22278
rect 15680 21242 15736 21244
rect 15760 21242 15816 21244
rect 15840 21242 15896 21244
rect 15920 21242 15976 21244
rect 15680 21190 15726 21242
rect 15726 21190 15736 21242
rect 15760 21190 15790 21242
rect 15790 21190 15802 21242
rect 15802 21190 15816 21242
rect 15840 21190 15854 21242
rect 15854 21190 15866 21242
rect 15866 21190 15896 21242
rect 15920 21190 15930 21242
rect 15930 21190 15976 21242
rect 15680 21188 15736 21190
rect 15760 21188 15816 21190
rect 15840 21188 15896 21190
rect 15920 21188 15976 21190
rect 15680 20154 15736 20156
rect 15760 20154 15816 20156
rect 15840 20154 15896 20156
rect 15920 20154 15976 20156
rect 15680 20102 15726 20154
rect 15726 20102 15736 20154
rect 15760 20102 15790 20154
rect 15790 20102 15802 20154
rect 15802 20102 15816 20154
rect 15840 20102 15854 20154
rect 15854 20102 15866 20154
rect 15866 20102 15896 20154
rect 15920 20102 15930 20154
rect 15930 20102 15976 20154
rect 15680 20100 15736 20102
rect 15760 20100 15816 20102
rect 15840 20100 15896 20102
rect 15920 20100 15976 20102
rect 15680 19066 15736 19068
rect 15760 19066 15816 19068
rect 15840 19066 15896 19068
rect 15920 19066 15976 19068
rect 15680 19014 15726 19066
rect 15726 19014 15736 19066
rect 15760 19014 15790 19066
rect 15790 19014 15802 19066
rect 15802 19014 15816 19066
rect 15840 19014 15854 19066
rect 15854 19014 15866 19066
rect 15866 19014 15896 19066
rect 15920 19014 15930 19066
rect 15930 19014 15976 19066
rect 15680 19012 15736 19014
rect 15760 19012 15816 19014
rect 15840 19012 15896 19014
rect 15920 19012 15976 19014
rect 15680 17978 15736 17980
rect 15760 17978 15816 17980
rect 15840 17978 15896 17980
rect 15920 17978 15976 17980
rect 15680 17926 15726 17978
rect 15726 17926 15736 17978
rect 15760 17926 15790 17978
rect 15790 17926 15802 17978
rect 15802 17926 15816 17978
rect 15840 17926 15854 17978
rect 15854 17926 15866 17978
rect 15866 17926 15896 17978
rect 15920 17926 15930 17978
rect 15930 17926 15976 17978
rect 15680 17924 15736 17926
rect 15760 17924 15816 17926
rect 15840 17924 15896 17926
rect 15920 17924 15976 17926
rect 15680 16890 15736 16892
rect 15760 16890 15816 16892
rect 15840 16890 15896 16892
rect 15920 16890 15976 16892
rect 15680 16838 15726 16890
rect 15726 16838 15736 16890
rect 15760 16838 15790 16890
rect 15790 16838 15802 16890
rect 15802 16838 15816 16890
rect 15840 16838 15854 16890
rect 15854 16838 15866 16890
rect 15866 16838 15896 16890
rect 15920 16838 15930 16890
rect 15930 16838 15976 16890
rect 15680 16836 15736 16838
rect 15760 16836 15816 16838
rect 15840 16836 15896 16838
rect 15920 16836 15976 16838
rect 15680 15802 15736 15804
rect 15760 15802 15816 15804
rect 15840 15802 15896 15804
rect 15920 15802 15976 15804
rect 15680 15750 15726 15802
rect 15726 15750 15736 15802
rect 15760 15750 15790 15802
rect 15790 15750 15802 15802
rect 15802 15750 15816 15802
rect 15840 15750 15854 15802
rect 15854 15750 15866 15802
rect 15866 15750 15896 15802
rect 15920 15750 15930 15802
rect 15930 15750 15976 15802
rect 15680 15748 15736 15750
rect 15760 15748 15816 15750
rect 15840 15748 15896 15750
rect 15920 15748 15976 15750
rect 15680 14714 15736 14716
rect 15760 14714 15816 14716
rect 15840 14714 15896 14716
rect 15920 14714 15976 14716
rect 15680 14662 15726 14714
rect 15726 14662 15736 14714
rect 15760 14662 15790 14714
rect 15790 14662 15802 14714
rect 15802 14662 15816 14714
rect 15840 14662 15854 14714
rect 15854 14662 15866 14714
rect 15866 14662 15896 14714
rect 15920 14662 15930 14714
rect 15930 14662 15976 14714
rect 15680 14660 15736 14662
rect 15760 14660 15816 14662
rect 15840 14660 15896 14662
rect 15920 14660 15976 14662
rect 15680 13626 15736 13628
rect 15760 13626 15816 13628
rect 15840 13626 15896 13628
rect 15920 13626 15976 13628
rect 15680 13574 15726 13626
rect 15726 13574 15736 13626
rect 15760 13574 15790 13626
rect 15790 13574 15802 13626
rect 15802 13574 15816 13626
rect 15840 13574 15854 13626
rect 15854 13574 15866 13626
rect 15866 13574 15896 13626
rect 15920 13574 15930 13626
rect 15930 13574 15976 13626
rect 15680 13572 15736 13574
rect 15760 13572 15816 13574
rect 15840 13572 15896 13574
rect 15920 13572 15976 13574
rect 15680 12538 15736 12540
rect 15760 12538 15816 12540
rect 15840 12538 15896 12540
rect 15920 12538 15976 12540
rect 15680 12486 15726 12538
rect 15726 12486 15736 12538
rect 15760 12486 15790 12538
rect 15790 12486 15802 12538
rect 15802 12486 15816 12538
rect 15840 12486 15854 12538
rect 15854 12486 15866 12538
rect 15866 12486 15896 12538
rect 15920 12486 15930 12538
rect 15930 12486 15976 12538
rect 15680 12484 15736 12486
rect 15760 12484 15816 12486
rect 15840 12484 15896 12486
rect 15920 12484 15976 12486
rect 15680 11450 15736 11452
rect 15760 11450 15816 11452
rect 15840 11450 15896 11452
rect 15920 11450 15976 11452
rect 15680 11398 15726 11450
rect 15726 11398 15736 11450
rect 15760 11398 15790 11450
rect 15790 11398 15802 11450
rect 15802 11398 15816 11450
rect 15840 11398 15854 11450
rect 15854 11398 15866 11450
rect 15866 11398 15896 11450
rect 15920 11398 15930 11450
rect 15930 11398 15976 11450
rect 15680 11396 15736 11398
rect 15760 11396 15816 11398
rect 15840 11396 15896 11398
rect 15920 11396 15976 11398
rect 15680 10362 15736 10364
rect 15760 10362 15816 10364
rect 15840 10362 15896 10364
rect 15920 10362 15976 10364
rect 15680 10310 15726 10362
rect 15726 10310 15736 10362
rect 15760 10310 15790 10362
rect 15790 10310 15802 10362
rect 15802 10310 15816 10362
rect 15840 10310 15854 10362
rect 15854 10310 15866 10362
rect 15866 10310 15896 10362
rect 15920 10310 15930 10362
rect 15930 10310 15976 10362
rect 15680 10308 15736 10310
rect 15760 10308 15816 10310
rect 15840 10308 15896 10310
rect 15920 10308 15976 10310
rect 15680 9274 15736 9276
rect 15760 9274 15816 9276
rect 15840 9274 15896 9276
rect 15920 9274 15976 9276
rect 15680 9222 15726 9274
rect 15726 9222 15736 9274
rect 15760 9222 15790 9274
rect 15790 9222 15802 9274
rect 15802 9222 15816 9274
rect 15840 9222 15854 9274
rect 15854 9222 15866 9274
rect 15866 9222 15896 9274
rect 15920 9222 15930 9274
rect 15930 9222 15976 9274
rect 15680 9220 15736 9222
rect 15760 9220 15816 9222
rect 15840 9220 15896 9222
rect 15920 9220 15976 9222
rect 15680 8186 15736 8188
rect 15760 8186 15816 8188
rect 15840 8186 15896 8188
rect 15920 8186 15976 8188
rect 15680 8134 15726 8186
rect 15726 8134 15736 8186
rect 15760 8134 15790 8186
rect 15790 8134 15802 8186
rect 15802 8134 15816 8186
rect 15840 8134 15854 8186
rect 15854 8134 15866 8186
rect 15866 8134 15896 8186
rect 15920 8134 15930 8186
rect 15930 8134 15976 8186
rect 15680 8132 15736 8134
rect 15760 8132 15816 8134
rect 15840 8132 15896 8134
rect 15920 8132 15976 8134
rect 15680 7098 15736 7100
rect 15760 7098 15816 7100
rect 15840 7098 15896 7100
rect 15920 7098 15976 7100
rect 15680 7046 15726 7098
rect 15726 7046 15736 7098
rect 15760 7046 15790 7098
rect 15790 7046 15802 7098
rect 15802 7046 15816 7098
rect 15840 7046 15854 7098
rect 15854 7046 15866 7098
rect 15866 7046 15896 7098
rect 15920 7046 15930 7098
rect 15930 7046 15976 7098
rect 15680 7044 15736 7046
rect 15760 7044 15816 7046
rect 15840 7044 15896 7046
rect 15920 7044 15976 7046
rect 15680 6010 15736 6012
rect 15760 6010 15816 6012
rect 15840 6010 15896 6012
rect 15920 6010 15976 6012
rect 15680 5958 15726 6010
rect 15726 5958 15736 6010
rect 15760 5958 15790 6010
rect 15790 5958 15802 6010
rect 15802 5958 15816 6010
rect 15840 5958 15854 6010
rect 15854 5958 15866 6010
rect 15866 5958 15896 6010
rect 15920 5958 15930 6010
rect 15930 5958 15976 6010
rect 15680 5956 15736 5958
rect 15760 5956 15816 5958
rect 15840 5956 15896 5958
rect 15920 5956 15976 5958
rect 15680 4922 15736 4924
rect 15760 4922 15816 4924
rect 15840 4922 15896 4924
rect 15920 4922 15976 4924
rect 15680 4870 15726 4922
rect 15726 4870 15736 4922
rect 15760 4870 15790 4922
rect 15790 4870 15802 4922
rect 15802 4870 15816 4922
rect 15840 4870 15854 4922
rect 15854 4870 15866 4922
rect 15866 4870 15896 4922
rect 15920 4870 15930 4922
rect 15930 4870 15976 4922
rect 15680 4868 15736 4870
rect 15760 4868 15816 4870
rect 15840 4868 15896 4870
rect 15920 4868 15976 4870
rect 15680 3834 15736 3836
rect 15760 3834 15816 3836
rect 15840 3834 15896 3836
rect 15920 3834 15976 3836
rect 15680 3782 15726 3834
rect 15726 3782 15736 3834
rect 15760 3782 15790 3834
rect 15790 3782 15802 3834
rect 15802 3782 15816 3834
rect 15840 3782 15854 3834
rect 15854 3782 15866 3834
rect 15866 3782 15896 3834
rect 15920 3782 15930 3834
rect 15930 3782 15976 3834
rect 15680 3780 15736 3782
rect 15760 3780 15816 3782
rect 15840 3780 15896 3782
rect 15920 3780 15976 3782
rect 15680 2746 15736 2748
rect 15760 2746 15816 2748
rect 15840 2746 15896 2748
rect 15920 2746 15976 2748
rect 15680 2694 15726 2746
rect 15726 2694 15736 2746
rect 15760 2694 15790 2746
rect 15790 2694 15802 2746
rect 15802 2694 15816 2746
rect 15840 2694 15854 2746
rect 15854 2694 15866 2746
rect 15866 2694 15896 2746
rect 15920 2694 15930 2746
rect 15930 2694 15976 2746
rect 15680 2692 15736 2694
rect 15760 2692 15816 2694
rect 15840 2692 15896 2694
rect 15920 2692 15976 2694
rect 16854 2488 16910 2544
rect 21178 27648 21234 27704
rect 19706 26696 19762 26752
rect 20626 27276 20628 27296
rect 20628 27276 20680 27296
rect 20680 27276 20682 27296
rect 20626 27240 20682 27276
rect 20718 26832 20774 26888
rect 23662 27512 23718 27568
rect 21914 27104 21970 27160
rect 21914 26968 21970 27024
rect 23570 27376 23626 27432
rect 25134 27104 25190 27160
rect 22466 26968 22522 27024
rect 26790 27004 26792 27024
rect 26792 27004 26844 27024
rect 26844 27004 26846 27024
rect 26790 26968 26846 27004
rect 22374 26696 22430 26752
rect 24122 26696 24178 26752
rect 22466 26560 22522 26616
rect 20350 26424 20406 26480
rect 22374 26324 22376 26344
rect 22376 26324 22428 26344
rect 22428 26324 22430 26344
rect 22374 26288 22430 26324
rect 24490 26308 24546 26344
rect 24490 26288 24492 26308
rect 24492 26288 24544 26308
rect 24544 26288 24546 26308
rect 29274 27784 29330 27840
rect 27158 26732 27160 26752
rect 27160 26732 27212 26752
rect 27212 26732 27214 26752
rect 27158 26696 27214 26732
rect 28170 26444 28226 26480
rect 28170 26424 28172 26444
rect 28172 26424 28224 26444
rect 28224 26424 28226 26444
rect 28998 26424 29054 26480
rect 29274 26732 29276 26752
rect 29276 26732 29328 26752
rect 29328 26732 29330 26752
rect 29274 26696 29330 26732
rect 30470 27376 30526 27432
rect 30654 27376 30710 27432
rect 30102 27240 30158 27296
rect 30194 27104 30250 27160
rect 30404 27226 30460 27228
rect 30484 27226 30540 27228
rect 30564 27226 30620 27228
rect 30644 27226 30700 27228
rect 30404 27174 30450 27226
rect 30450 27174 30460 27226
rect 30484 27174 30514 27226
rect 30514 27174 30526 27226
rect 30526 27174 30540 27226
rect 30564 27174 30578 27226
rect 30578 27174 30590 27226
rect 30590 27174 30620 27226
rect 30644 27174 30654 27226
rect 30654 27174 30700 27226
rect 30404 27172 30460 27174
rect 30484 27172 30540 27174
rect 30564 27172 30620 27174
rect 30644 27172 30700 27174
rect 31114 27532 31170 27568
rect 31114 27512 31116 27532
rect 31116 27512 31168 27532
rect 31168 27512 31170 27532
rect 31390 27548 31392 27568
rect 31392 27548 31444 27568
rect 31444 27548 31446 27568
rect 31390 27512 31446 27548
rect 17314 1536 17370 1592
rect 19706 2372 19762 2408
rect 19706 2352 19708 2372
rect 19708 2352 19760 2372
rect 19760 2352 19762 2372
rect 26146 1672 26202 1728
rect 28170 2352 28226 2408
rect 30404 26138 30460 26140
rect 30484 26138 30540 26140
rect 30564 26138 30620 26140
rect 30644 26138 30700 26140
rect 30404 26086 30450 26138
rect 30450 26086 30460 26138
rect 30484 26086 30514 26138
rect 30514 26086 30526 26138
rect 30526 26086 30540 26138
rect 30564 26086 30578 26138
rect 30578 26086 30590 26138
rect 30590 26086 30620 26138
rect 30644 26086 30654 26138
rect 30654 26086 30700 26138
rect 30404 26084 30460 26086
rect 30484 26084 30540 26086
rect 30564 26084 30620 26086
rect 30644 26084 30700 26086
rect 30404 25050 30460 25052
rect 30484 25050 30540 25052
rect 30564 25050 30620 25052
rect 30644 25050 30700 25052
rect 30404 24998 30450 25050
rect 30450 24998 30460 25050
rect 30484 24998 30514 25050
rect 30514 24998 30526 25050
rect 30526 24998 30540 25050
rect 30564 24998 30578 25050
rect 30578 24998 30590 25050
rect 30590 24998 30620 25050
rect 30644 24998 30654 25050
rect 30654 24998 30700 25050
rect 30404 24996 30460 24998
rect 30484 24996 30540 24998
rect 30564 24996 30620 24998
rect 30644 24996 30700 24998
rect 30404 23962 30460 23964
rect 30484 23962 30540 23964
rect 30564 23962 30620 23964
rect 30644 23962 30700 23964
rect 30404 23910 30450 23962
rect 30450 23910 30460 23962
rect 30484 23910 30514 23962
rect 30514 23910 30526 23962
rect 30526 23910 30540 23962
rect 30564 23910 30578 23962
rect 30578 23910 30590 23962
rect 30590 23910 30620 23962
rect 30644 23910 30654 23962
rect 30654 23910 30700 23962
rect 30404 23908 30460 23910
rect 30484 23908 30540 23910
rect 30564 23908 30620 23910
rect 30644 23908 30700 23910
rect 30404 22874 30460 22876
rect 30484 22874 30540 22876
rect 30564 22874 30620 22876
rect 30644 22874 30700 22876
rect 30404 22822 30450 22874
rect 30450 22822 30460 22874
rect 30484 22822 30514 22874
rect 30514 22822 30526 22874
rect 30526 22822 30540 22874
rect 30564 22822 30578 22874
rect 30578 22822 30590 22874
rect 30590 22822 30620 22874
rect 30644 22822 30654 22874
rect 30654 22822 30700 22874
rect 30404 22820 30460 22822
rect 30484 22820 30540 22822
rect 30564 22820 30620 22822
rect 30644 22820 30700 22822
rect 32126 27396 32182 27432
rect 32126 27376 32128 27396
rect 32128 27376 32180 27396
rect 32180 27376 32182 27396
rect 31574 26968 31630 27024
rect 30404 21786 30460 21788
rect 30484 21786 30540 21788
rect 30564 21786 30620 21788
rect 30644 21786 30700 21788
rect 30404 21734 30450 21786
rect 30450 21734 30460 21786
rect 30484 21734 30514 21786
rect 30514 21734 30526 21786
rect 30526 21734 30540 21786
rect 30564 21734 30578 21786
rect 30578 21734 30590 21786
rect 30590 21734 30620 21786
rect 30644 21734 30654 21786
rect 30654 21734 30700 21786
rect 30404 21732 30460 21734
rect 30484 21732 30540 21734
rect 30564 21732 30620 21734
rect 30644 21732 30700 21734
rect 30404 20698 30460 20700
rect 30484 20698 30540 20700
rect 30564 20698 30620 20700
rect 30644 20698 30700 20700
rect 30404 20646 30450 20698
rect 30450 20646 30460 20698
rect 30484 20646 30514 20698
rect 30514 20646 30526 20698
rect 30526 20646 30540 20698
rect 30564 20646 30578 20698
rect 30578 20646 30590 20698
rect 30590 20646 30620 20698
rect 30644 20646 30654 20698
rect 30654 20646 30700 20698
rect 30404 20644 30460 20646
rect 30484 20644 30540 20646
rect 30564 20644 30620 20646
rect 30644 20644 30700 20646
rect 30404 19610 30460 19612
rect 30484 19610 30540 19612
rect 30564 19610 30620 19612
rect 30644 19610 30700 19612
rect 30404 19558 30450 19610
rect 30450 19558 30460 19610
rect 30484 19558 30514 19610
rect 30514 19558 30526 19610
rect 30526 19558 30540 19610
rect 30564 19558 30578 19610
rect 30578 19558 30590 19610
rect 30590 19558 30620 19610
rect 30644 19558 30654 19610
rect 30654 19558 30700 19610
rect 30404 19556 30460 19558
rect 30484 19556 30540 19558
rect 30564 19556 30620 19558
rect 30644 19556 30700 19558
rect 30404 18522 30460 18524
rect 30484 18522 30540 18524
rect 30564 18522 30620 18524
rect 30644 18522 30700 18524
rect 30404 18470 30450 18522
rect 30450 18470 30460 18522
rect 30484 18470 30514 18522
rect 30514 18470 30526 18522
rect 30526 18470 30540 18522
rect 30564 18470 30578 18522
rect 30578 18470 30590 18522
rect 30590 18470 30620 18522
rect 30644 18470 30654 18522
rect 30654 18470 30700 18522
rect 30404 18468 30460 18470
rect 30484 18468 30540 18470
rect 30564 18468 30620 18470
rect 30644 18468 30700 18470
rect 30404 17434 30460 17436
rect 30484 17434 30540 17436
rect 30564 17434 30620 17436
rect 30644 17434 30700 17436
rect 30404 17382 30450 17434
rect 30450 17382 30460 17434
rect 30484 17382 30514 17434
rect 30514 17382 30526 17434
rect 30526 17382 30540 17434
rect 30564 17382 30578 17434
rect 30578 17382 30590 17434
rect 30590 17382 30620 17434
rect 30644 17382 30654 17434
rect 30654 17382 30700 17434
rect 30404 17380 30460 17382
rect 30484 17380 30540 17382
rect 30564 17380 30620 17382
rect 30644 17380 30700 17382
rect 30404 16346 30460 16348
rect 30484 16346 30540 16348
rect 30564 16346 30620 16348
rect 30644 16346 30700 16348
rect 30404 16294 30450 16346
rect 30450 16294 30460 16346
rect 30484 16294 30514 16346
rect 30514 16294 30526 16346
rect 30526 16294 30540 16346
rect 30564 16294 30578 16346
rect 30578 16294 30590 16346
rect 30590 16294 30620 16346
rect 30644 16294 30654 16346
rect 30654 16294 30700 16346
rect 30404 16292 30460 16294
rect 30484 16292 30540 16294
rect 30564 16292 30620 16294
rect 30644 16292 30700 16294
rect 30404 15258 30460 15260
rect 30484 15258 30540 15260
rect 30564 15258 30620 15260
rect 30644 15258 30700 15260
rect 30404 15206 30450 15258
rect 30450 15206 30460 15258
rect 30484 15206 30514 15258
rect 30514 15206 30526 15258
rect 30526 15206 30540 15258
rect 30564 15206 30578 15258
rect 30578 15206 30590 15258
rect 30590 15206 30620 15258
rect 30644 15206 30654 15258
rect 30654 15206 30700 15258
rect 30404 15204 30460 15206
rect 30484 15204 30540 15206
rect 30564 15204 30620 15206
rect 30644 15204 30700 15206
rect 30404 14170 30460 14172
rect 30484 14170 30540 14172
rect 30564 14170 30620 14172
rect 30644 14170 30700 14172
rect 30404 14118 30450 14170
rect 30450 14118 30460 14170
rect 30484 14118 30514 14170
rect 30514 14118 30526 14170
rect 30526 14118 30540 14170
rect 30564 14118 30578 14170
rect 30578 14118 30590 14170
rect 30590 14118 30620 14170
rect 30644 14118 30654 14170
rect 30654 14118 30700 14170
rect 30404 14116 30460 14118
rect 30484 14116 30540 14118
rect 30564 14116 30620 14118
rect 30644 14116 30700 14118
rect 30404 13082 30460 13084
rect 30484 13082 30540 13084
rect 30564 13082 30620 13084
rect 30644 13082 30700 13084
rect 30404 13030 30450 13082
rect 30450 13030 30460 13082
rect 30484 13030 30514 13082
rect 30514 13030 30526 13082
rect 30526 13030 30540 13082
rect 30564 13030 30578 13082
rect 30578 13030 30590 13082
rect 30590 13030 30620 13082
rect 30644 13030 30654 13082
rect 30654 13030 30700 13082
rect 30404 13028 30460 13030
rect 30484 13028 30540 13030
rect 30564 13028 30620 13030
rect 30644 13028 30700 13030
rect 30404 11994 30460 11996
rect 30484 11994 30540 11996
rect 30564 11994 30620 11996
rect 30644 11994 30700 11996
rect 30404 11942 30450 11994
rect 30450 11942 30460 11994
rect 30484 11942 30514 11994
rect 30514 11942 30526 11994
rect 30526 11942 30540 11994
rect 30564 11942 30578 11994
rect 30578 11942 30590 11994
rect 30590 11942 30620 11994
rect 30644 11942 30654 11994
rect 30654 11942 30700 11994
rect 30404 11940 30460 11942
rect 30484 11940 30540 11942
rect 30564 11940 30620 11942
rect 30644 11940 30700 11942
rect 30404 10906 30460 10908
rect 30484 10906 30540 10908
rect 30564 10906 30620 10908
rect 30644 10906 30700 10908
rect 30404 10854 30450 10906
rect 30450 10854 30460 10906
rect 30484 10854 30514 10906
rect 30514 10854 30526 10906
rect 30526 10854 30540 10906
rect 30564 10854 30578 10906
rect 30578 10854 30590 10906
rect 30590 10854 30620 10906
rect 30644 10854 30654 10906
rect 30654 10854 30700 10906
rect 30404 10852 30460 10854
rect 30484 10852 30540 10854
rect 30564 10852 30620 10854
rect 30644 10852 30700 10854
rect 31482 26580 31538 26616
rect 31482 26560 31484 26580
rect 31484 26560 31536 26580
rect 31536 26560 31538 26580
rect 31574 26288 31630 26344
rect 31850 26288 31906 26344
rect 32034 26288 32090 26344
rect 30404 9818 30460 9820
rect 30484 9818 30540 9820
rect 30564 9818 30620 9820
rect 30644 9818 30700 9820
rect 30404 9766 30450 9818
rect 30450 9766 30460 9818
rect 30484 9766 30514 9818
rect 30514 9766 30526 9818
rect 30526 9766 30540 9818
rect 30564 9766 30578 9818
rect 30578 9766 30590 9818
rect 30590 9766 30620 9818
rect 30644 9766 30654 9818
rect 30654 9766 30700 9818
rect 30404 9764 30460 9766
rect 30484 9764 30540 9766
rect 30564 9764 30620 9766
rect 30644 9764 30700 9766
rect 30404 8730 30460 8732
rect 30484 8730 30540 8732
rect 30564 8730 30620 8732
rect 30644 8730 30700 8732
rect 30404 8678 30450 8730
rect 30450 8678 30460 8730
rect 30484 8678 30514 8730
rect 30514 8678 30526 8730
rect 30526 8678 30540 8730
rect 30564 8678 30578 8730
rect 30578 8678 30590 8730
rect 30590 8678 30620 8730
rect 30644 8678 30654 8730
rect 30654 8678 30700 8730
rect 30404 8676 30460 8678
rect 30484 8676 30540 8678
rect 30564 8676 30620 8678
rect 30644 8676 30700 8678
rect 30404 7642 30460 7644
rect 30484 7642 30540 7644
rect 30564 7642 30620 7644
rect 30644 7642 30700 7644
rect 30404 7590 30450 7642
rect 30450 7590 30460 7642
rect 30484 7590 30514 7642
rect 30514 7590 30526 7642
rect 30526 7590 30540 7642
rect 30564 7590 30578 7642
rect 30578 7590 30590 7642
rect 30590 7590 30620 7642
rect 30644 7590 30654 7642
rect 30654 7590 30700 7642
rect 30404 7588 30460 7590
rect 30484 7588 30540 7590
rect 30564 7588 30620 7590
rect 30644 7588 30700 7590
rect 30404 6554 30460 6556
rect 30484 6554 30540 6556
rect 30564 6554 30620 6556
rect 30644 6554 30700 6556
rect 30404 6502 30450 6554
rect 30450 6502 30460 6554
rect 30484 6502 30514 6554
rect 30514 6502 30526 6554
rect 30526 6502 30540 6554
rect 30564 6502 30578 6554
rect 30578 6502 30590 6554
rect 30590 6502 30620 6554
rect 30644 6502 30654 6554
rect 30654 6502 30700 6554
rect 30404 6500 30460 6502
rect 30484 6500 30540 6502
rect 30564 6500 30620 6502
rect 30644 6500 30700 6502
rect 30404 5466 30460 5468
rect 30484 5466 30540 5468
rect 30564 5466 30620 5468
rect 30644 5466 30700 5468
rect 30404 5414 30450 5466
rect 30450 5414 30460 5466
rect 30484 5414 30514 5466
rect 30514 5414 30526 5466
rect 30526 5414 30540 5466
rect 30564 5414 30578 5466
rect 30578 5414 30590 5466
rect 30590 5414 30620 5466
rect 30644 5414 30654 5466
rect 30654 5414 30700 5466
rect 30404 5412 30460 5414
rect 30484 5412 30540 5414
rect 30564 5412 30620 5414
rect 30644 5412 30700 5414
rect 30404 4378 30460 4380
rect 30484 4378 30540 4380
rect 30564 4378 30620 4380
rect 30644 4378 30700 4380
rect 30404 4326 30450 4378
rect 30450 4326 30460 4378
rect 30484 4326 30514 4378
rect 30514 4326 30526 4378
rect 30526 4326 30540 4378
rect 30564 4326 30578 4378
rect 30578 4326 30590 4378
rect 30590 4326 30620 4378
rect 30644 4326 30654 4378
rect 30654 4326 30700 4378
rect 30404 4324 30460 4326
rect 30484 4324 30540 4326
rect 30564 4324 30620 4326
rect 30644 4324 30700 4326
rect 33046 27548 33048 27568
rect 33048 27548 33100 27568
rect 33100 27548 33102 27568
rect 33046 27512 33102 27548
rect 34058 27648 34114 27704
rect 33598 27240 33654 27296
rect 33598 26560 33654 26616
rect 34610 26988 34666 27024
rect 34610 26968 34612 26988
rect 34612 26968 34664 26988
rect 34664 26968 34666 26988
rect 33874 26424 33930 26480
rect 34978 26560 35034 26616
rect 35346 27376 35402 27432
rect 35254 26968 35310 27024
rect 35162 26560 35218 26616
rect 37922 27396 37978 27432
rect 37922 27376 37924 27396
rect 37924 27376 37976 27396
rect 37976 27376 37978 27396
rect 35806 26444 35862 26480
rect 35806 26424 35808 26444
rect 35808 26424 35860 26444
rect 35860 26424 35862 26444
rect 38290 27784 38346 27840
rect 38382 26560 38438 26616
rect 30404 3290 30460 3292
rect 30484 3290 30540 3292
rect 30564 3290 30620 3292
rect 30644 3290 30700 3292
rect 30404 3238 30450 3290
rect 30450 3238 30460 3290
rect 30484 3238 30514 3290
rect 30514 3238 30526 3290
rect 30526 3238 30540 3290
rect 30564 3238 30578 3290
rect 30578 3238 30590 3290
rect 30590 3238 30620 3290
rect 30644 3238 30654 3290
rect 30654 3238 30700 3290
rect 30404 3236 30460 3238
rect 30484 3236 30540 3238
rect 30564 3236 30620 3238
rect 30644 3236 30700 3238
rect 28446 1536 28502 1592
rect 30404 2202 30460 2204
rect 30484 2202 30540 2204
rect 30564 2202 30620 2204
rect 30644 2202 30700 2204
rect 30404 2150 30450 2202
rect 30450 2150 30460 2202
rect 30484 2150 30514 2202
rect 30514 2150 30526 2202
rect 30526 2150 30540 2202
rect 30564 2150 30578 2202
rect 30578 2150 30590 2202
rect 30590 2150 30620 2202
rect 30644 2150 30654 2202
rect 30654 2150 30700 2202
rect 30404 2148 30460 2150
rect 30484 2148 30540 2150
rect 30564 2148 30620 2150
rect 30644 2148 30700 2150
rect 30746 1808 30802 1864
rect 1398 720 1454 776
rect 31574 1672 31630 1728
rect 40222 27920 40278 27976
rect 38566 26424 38622 26480
rect 40682 27548 40684 27568
rect 40684 27548 40736 27568
rect 40736 27548 40738 27568
rect 40682 27512 40738 27548
rect 40314 27124 40370 27160
rect 40314 27104 40316 27124
rect 40316 27104 40368 27124
rect 40368 27104 40370 27124
rect 40774 26016 40830 26072
rect 40038 3032 40094 3088
rect 38566 1808 38622 1864
rect 39854 2896 39910 2952
rect 39578 2352 39634 2408
rect 40314 3576 40370 3632
rect 43810 27532 43866 27568
rect 43810 27512 43812 27532
rect 43812 27512 43864 27532
rect 43864 27512 43866 27532
rect 45128 27770 45184 27772
rect 45208 27770 45264 27772
rect 45288 27770 45344 27772
rect 45368 27770 45424 27772
rect 45128 27718 45174 27770
rect 45174 27718 45184 27770
rect 45208 27718 45238 27770
rect 45238 27718 45250 27770
rect 45250 27718 45264 27770
rect 45288 27718 45302 27770
rect 45302 27718 45314 27770
rect 45314 27718 45344 27770
rect 45368 27718 45378 27770
rect 45378 27718 45424 27770
rect 45128 27716 45184 27718
rect 45208 27716 45264 27718
rect 45288 27716 45344 27718
rect 45368 27716 45424 27718
rect 41878 27104 41934 27160
rect 40958 26696 41014 26752
rect 41142 26560 41198 26616
rect 40958 26424 41014 26480
rect 41234 26288 41290 26344
rect 41786 26288 41842 26344
rect 41234 3188 41290 3224
rect 41234 3168 41236 3188
rect 41236 3168 41288 3188
rect 41288 3168 41290 3188
rect 45926 27104 45982 27160
rect 45128 26682 45184 26684
rect 45208 26682 45264 26684
rect 45288 26682 45344 26684
rect 45368 26682 45424 26684
rect 45128 26630 45174 26682
rect 45174 26630 45184 26682
rect 45208 26630 45238 26682
rect 45238 26630 45250 26682
rect 45250 26630 45264 26682
rect 45288 26630 45302 26682
rect 45302 26630 45314 26682
rect 45314 26630 45344 26682
rect 45368 26630 45378 26682
rect 45378 26630 45424 26682
rect 45128 26628 45184 26630
rect 45208 26628 45264 26630
rect 45288 26628 45344 26630
rect 45368 26628 45424 26630
rect 44086 26560 44142 26616
rect 43442 26460 43444 26480
rect 43444 26460 43496 26480
rect 43496 26460 43498 26480
rect 43442 26424 43498 26460
rect 49054 27784 49110 27840
rect 45128 25594 45184 25596
rect 45208 25594 45264 25596
rect 45288 25594 45344 25596
rect 45368 25594 45424 25596
rect 45128 25542 45174 25594
rect 45174 25542 45184 25594
rect 45208 25542 45238 25594
rect 45238 25542 45250 25594
rect 45250 25542 45264 25594
rect 45288 25542 45302 25594
rect 45302 25542 45314 25594
rect 45314 25542 45344 25594
rect 45368 25542 45378 25594
rect 45378 25542 45424 25594
rect 45128 25540 45184 25542
rect 45208 25540 45264 25542
rect 45288 25540 45344 25542
rect 45368 25540 45424 25542
rect 45128 24506 45184 24508
rect 45208 24506 45264 24508
rect 45288 24506 45344 24508
rect 45368 24506 45424 24508
rect 45128 24454 45174 24506
rect 45174 24454 45184 24506
rect 45208 24454 45238 24506
rect 45238 24454 45250 24506
rect 45250 24454 45264 24506
rect 45288 24454 45302 24506
rect 45302 24454 45314 24506
rect 45314 24454 45344 24506
rect 45368 24454 45378 24506
rect 45378 24454 45424 24506
rect 45128 24452 45184 24454
rect 45208 24452 45264 24454
rect 45288 24452 45344 24454
rect 45368 24452 45424 24454
rect 45128 23418 45184 23420
rect 45208 23418 45264 23420
rect 45288 23418 45344 23420
rect 45368 23418 45424 23420
rect 45128 23366 45174 23418
rect 45174 23366 45184 23418
rect 45208 23366 45238 23418
rect 45238 23366 45250 23418
rect 45250 23366 45264 23418
rect 45288 23366 45302 23418
rect 45302 23366 45314 23418
rect 45314 23366 45344 23418
rect 45368 23366 45378 23418
rect 45378 23366 45424 23418
rect 45128 23364 45184 23366
rect 45208 23364 45264 23366
rect 45288 23364 45344 23366
rect 45368 23364 45424 23366
rect 45128 22330 45184 22332
rect 45208 22330 45264 22332
rect 45288 22330 45344 22332
rect 45368 22330 45424 22332
rect 45128 22278 45174 22330
rect 45174 22278 45184 22330
rect 45208 22278 45238 22330
rect 45238 22278 45250 22330
rect 45250 22278 45264 22330
rect 45288 22278 45302 22330
rect 45302 22278 45314 22330
rect 45314 22278 45344 22330
rect 45368 22278 45378 22330
rect 45378 22278 45424 22330
rect 45128 22276 45184 22278
rect 45208 22276 45264 22278
rect 45288 22276 45344 22278
rect 45368 22276 45424 22278
rect 45128 21242 45184 21244
rect 45208 21242 45264 21244
rect 45288 21242 45344 21244
rect 45368 21242 45424 21244
rect 45128 21190 45174 21242
rect 45174 21190 45184 21242
rect 45208 21190 45238 21242
rect 45238 21190 45250 21242
rect 45250 21190 45264 21242
rect 45288 21190 45302 21242
rect 45302 21190 45314 21242
rect 45314 21190 45344 21242
rect 45368 21190 45378 21242
rect 45378 21190 45424 21242
rect 45128 21188 45184 21190
rect 45208 21188 45264 21190
rect 45288 21188 45344 21190
rect 45368 21188 45424 21190
rect 45128 20154 45184 20156
rect 45208 20154 45264 20156
rect 45288 20154 45344 20156
rect 45368 20154 45424 20156
rect 45128 20102 45174 20154
rect 45174 20102 45184 20154
rect 45208 20102 45238 20154
rect 45238 20102 45250 20154
rect 45250 20102 45264 20154
rect 45288 20102 45302 20154
rect 45302 20102 45314 20154
rect 45314 20102 45344 20154
rect 45368 20102 45378 20154
rect 45378 20102 45424 20154
rect 45128 20100 45184 20102
rect 45208 20100 45264 20102
rect 45288 20100 45344 20102
rect 45368 20100 45424 20102
rect 45128 19066 45184 19068
rect 45208 19066 45264 19068
rect 45288 19066 45344 19068
rect 45368 19066 45424 19068
rect 45128 19014 45174 19066
rect 45174 19014 45184 19066
rect 45208 19014 45238 19066
rect 45238 19014 45250 19066
rect 45250 19014 45264 19066
rect 45288 19014 45302 19066
rect 45302 19014 45314 19066
rect 45314 19014 45344 19066
rect 45368 19014 45378 19066
rect 45378 19014 45424 19066
rect 45128 19012 45184 19014
rect 45208 19012 45264 19014
rect 45288 19012 45344 19014
rect 45368 19012 45424 19014
rect 45128 17978 45184 17980
rect 45208 17978 45264 17980
rect 45288 17978 45344 17980
rect 45368 17978 45424 17980
rect 45128 17926 45174 17978
rect 45174 17926 45184 17978
rect 45208 17926 45238 17978
rect 45238 17926 45250 17978
rect 45250 17926 45264 17978
rect 45288 17926 45302 17978
rect 45302 17926 45314 17978
rect 45314 17926 45344 17978
rect 45368 17926 45378 17978
rect 45378 17926 45424 17978
rect 45128 17924 45184 17926
rect 45208 17924 45264 17926
rect 45288 17924 45344 17926
rect 45368 17924 45424 17926
rect 45128 16890 45184 16892
rect 45208 16890 45264 16892
rect 45288 16890 45344 16892
rect 45368 16890 45424 16892
rect 45128 16838 45174 16890
rect 45174 16838 45184 16890
rect 45208 16838 45238 16890
rect 45238 16838 45250 16890
rect 45250 16838 45264 16890
rect 45288 16838 45302 16890
rect 45302 16838 45314 16890
rect 45314 16838 45344 16890
rect 45368 16838 45378 16890
rect 45378 16838 45424 16890
rect 45128 16836 45184 16838
rect 45208 16836 45264 16838
rect 45288 16836 45344 16838
rect 45368 16836 45424 16838
rect 45128 15802 45184 15804
rect 45208 15802 45264 15804
rect 45288 15802 45344 15804
rect 45368 15802 45424 15804
rect 45128 15750 45174 15802
rect 45174 15750 45184 15802
rect 45208 15750 45238 15802
rect 45238 15750 45250 15802
rect 45250 15750 45264 15802
rect 45288 15750 45302 15802
rect 45302 15750 45314 15802
rect 45314 15750 45344 15802
rect 45368 15750 45378 15802
rect 45378 15750 45424 15802
rect 45128 15748 45184 15750
rect 45208 15748 45264 15750
rect 45288 15748 45344 15750
rect 45368 15748 45424 15750
rect 45128 14714 45184 14716
rect 45208 14714 45264 14716
rect 45288 14714 45344 14716
rect 45368 14714 45424 14716
rect 45128 14662 45174 14714
rect 45174 14662 45184 14714
rect 45208 14662 45238 14714
rect 45238 14662 45250 14714
rect 45250 14662 45264 14714
rect 45288 14662 45302 14714
rect 45302 14662 45314 14714
rect 45314 14662 45344 14714
rect 45368 14662 45378 14714
rect 45378 14662 45424 14714
rect 45128 14660 45184 14662
rect 45208 14660 45264 14662
rect 45288 14660 45344 14662
rect 45368 14660 45424 14662
rect 45128 13626 45184 13628
rect 45208 13626 45264 13628
rect 45288 13626 45344 13628
rect 45368 13626 45424 13628
rect 45128 13574 45174 13626
rect 45174 13574 45184 13626
rect 45208 13574 45238 13626
rect 45238 13574 45250 13626
rect 45250 13574 45264 13626
rect 45288 13574 45302 13626
rect 45302 13574 45314 13626
rect 45314 13574 45344 13626
rect 45368 13574 45378 13626
rect 45378 13574 45424 13626
rect 45128 13572 45184 13574
rect 45208 13572 45264 13574
rect 45288 13572 45344 13574
rect 45368 13572 45424 13574
rect 42430 3476 42432 3496
rect 42432 3476 42484 3496
rect 42484 3476 42486 3496
rect 42430 3440 42486 3476
rect 45128 12538 45184 12540
rect 45208 12538 45264 12540
rect 45288 12538 45344 12540
rect 45368 12538 45424 12540
rect 45128 12486 45174 12538
rect 45174 12486 45184 12538
rect 45208 12486 45238 12538
rect 45238 12486 45250 12538
rect 45250 12486 45264 12538
rect 45288 12486 45302 12538
rect 45302 12486 45314 12538
rect 45314 12486 45344 12538
rect 45368 12486 45378 12538
rect 45378 12486 45424 12538
rect 45128 12484 45184 12486
rect 45208 12484 45264 12486
rect 45288 12484 45344 12486
rect 45368 12484 45424 12486
rect 45128 11450 45184 11452
rect 45208 11450 45264 11452
rect 45288 11450 45344 11452
rect 45368 11450 45424 11452
rect 45128 11398 45174 11450
rect 45174 11398 45184 11450
rect 45208 11398 45238 11450
rect 45238 11398 45250 11450
rect 45250 11398 45264 11450
rect 45288 11398 45302 11450
rect 45302 11398 45314 11450
rect 45314 11398 45344 11450
rect 45368 11398 45378 11450
rect 45378 11398 45424 11450
rect 45128 11396 45184 11398
rect 45208 11396 45264 11398
rect 45288 11396 45344 11398
rect 45368 11396 45424 11398
rect 45128 10362 45184 10364
rect 45208 10362 45264 10364
rect 45288 10362 45344 10364
rect 45368 10362 45424 10364
rect 45128 10310 45174 10362
rect 45174 10310 45184 10362
rect 45208 10310 45238 10362
rect 45238 10310 45250 10362
rect 45250 10310 45264 10362
rect 45288 10310 45302 10362
rect 45302 10310 45314 10362
rect 45314 10310 45344 10362
rect 45368 10310 45378 10362
rect 45378 10310 45424 10362
rect 45128 10308 45184 10310
rect 45208 10308 45264 10310
rect 45288 10308 45344 10310
rect 45368 10308 45424 10310
rect 45128 9274 45184 9276
rect 45208 9274 45264 9276
rect 45288 9274 45344 9276
rect 45368 9274 45424 9276
rect 45128 9222 45174 9274
rect 45174 9222 45184 9274
rect 45208 9222 45238 9274
rect 45238 9222 45250 9274
rect 45250 9222 45264 9274
rect 45288 9222 45302 9274
rect 45302 9222 45314 9274
rect 45314 9222 45344 9274
rect 45368 9222 45378 9274
rect 45378 9222 45424 9274
rect 45128 9220 45184 9222
rect 45208 9220 45264 9222
rect 45288 9220 45344 9222
rect 45368 9220 45424 9222
rect 45128 8186 45184 8188
rect 45208 8186 45264 8188
rect 45288 8186 45344 8188
rect 45368 8186 45424 8188
rect 45128 8134 45174 8186
rect 45174 8134 45184 8186
rect 45208 8134 45238 8186
rect 45238 8134 45250 8186
rect 45250 8134 45264 8186
rect 45288 8134 45302 8186
rect 45302 8134 45314 8186
rect 45314 8134 45344 8186
rect 45368 8134 45378 8186
rect 45378 8134 45424 8186
rect 45128 8132 45184 8134
rect 45208 8132 45264 8134
rect 45288 8132 45344 8134
rect 45368 8132 45424 8134
rect 47122 26152 47178 26208
rect 47306 26016 47362 26072
rect 45128 7098 45184 7100
rect 45208 7098 45264 7100
rect 45288 7098 45344 7100
rect 45368 7098 45424 7100
rect 45128 7046 45174 7098
rect 45174 7046 45184 7098
rect 45208 7046 45238 7098
rect 45238 7046 45250 7098
rect 45250 7046 45264 7098
rect 45288 7046 45302 7098
rect 45302 7046 45314 7098
rect 45314 7046 45344 7098
rect 45368 7046 45378 7098
rect 45378 7046 45424 7098
rect 45128 7044 45184 7046
rect 45208 7044 45264 7046
rect 45288 7044 45344 7046
rect 45368 7044 45424 7046
rect 45128 6010 45184 6012
rect 45208 6010 45264 6012
rect 45288 6010 45344 6012
rect 45368 6010 45424 6012
rect 45128 5958 45174 6010
rect 45174 5958 45184 6010
rect 45208 5958 45238 6010
rect 45238 5958 45250 6010
rect 45250 5958 45264 6010
rect 45288 5958 45302 6010
rect 45302 5958 45314 6010
rect 45314 5958 45344 6010
rect 45368 5958 45378 6010
rect 45378 5958 45424 6010
rect 45128 5956 45184 5958
rect 45208 5956 45264 5958
rect 45288 5956 45344 5958
rect 45368 5956 45424 5958
rect 45128 4922 45184 4924
rect 45208 4922 45264 4924
rect 45288 4922 45344 4924
rect 45368 4922 45424 4924
rect 45128 4870 45174 4922
rect 45174 4870 45184 4922
rect 45208 4870 45238 4922
rect 45238 4870 45250 4922
rect 45250 4870 45264 4922
rect 45288 4870 45302 4922
rect 45302 4870 45314 4922
rect 45314 4870 45344 4922
rect 45368 4870 45378 4922
rect 45378 4870 45424 4922
rect 45128 4868 45184 4870
rect 45208 4868 45264 4870
rect 45288 4868 45344 4870
rect 45368 4868 45424 4870
rect 45128 3834 45184 3836
rect 45208 3834 45264 3836
rect 45288 3834 45344 3836
rect 45368 3834 45424 3836
rect 45128 3782 45174 3834
rect 45174 3782 45184 3834
rect 45208 3782 45238 3834
rect 45238 3782 45250 3834
rect 45250 3782 45264 3834
rect 45288 3782 45302 3834
rect 45302 3782 45314 3834
rect 45314 3782 45344 3834
rect 45368 3782 45378 3834
rect 45378 3782 45424 3834
rect 45128 3780 45184 3782
rect 45208 3780 45264 3782
rect 45288 3780 45344 3782
rect 45368 3780 45424 3782
rect 43258 3304 43314 3360
rect 45374 3052 45430 3088
rect 45374 3032 45376 3052
rect 45376 3032 45428 3052
rect 45428 3032 45430 3052
rect 45128 2746 45184 2748
rect 45208 2746 45264 2748
rect 45288 2746 45344 2748
rect 45368 2746 45424 2748
rect 45128 2694 45174 2746
rect 45174 2694 45184 2746
rect 45208 2694 45238 2746
rect 45238 2694 45250 2746
rect 45250 2694 45264 2746
rect 45288 2694 45302 2746
rect 45302 2694 45314 2746
rect 45314 2694 45344 2746
rect 45368 2694 45378 2746
rect 45378 2694 45424 2746
rect 45128 2692 45184 2694
rect 45208 2692 45264 2694
rect 45288 2692 45344 2694
rect 45368 2692 45424 2694
rect 46202 3168 46258 3224
rect 47306 3576 47362 3632
rect 46754 2372 46810 2408
rect 46754 2352 46756 2372
rect 46756 2352 46808 2372
rect 46808 2352 46810 2372
rect 48042 3476 48044 3496
rect 48044 3476 48096 3496
rect 48096 3476 48098 3496
rect 47582 3340 47584 3360
rect 47584 3340 47636 3360
rect 47636 3340 47638 3360
rect 47582 3304 47638 3340
rect 48042 3440 48098 3476
rect 47490 2896 47546 2952
rect 47950 2352 48006 2408
rect 50250 27512 50306 27568
rect 50434 27512 50490 27568
rect 50158 26424 50214 26480
rect 50158 26288 50214 26344
rect 50434 27240 50490 27296
rect 50618 27240 50674 27296
rect 51814 27512 51870 27568
rect 50894 27104 50950 27160
rect 50618 26696 50674 26752
rect 50526 26560 50582 26616
rect 50710 26424 50766 26480
rect 50986 26308 51042 26344
rect 50986 26288 50988 26308
rect 50988 26288 51040 26308
rect 51040 26288 51042 26308
rect 50894 26152 50950 26208
rect 51170 26696 51226 26752
rect 51262 26560 51318 26616
rect 51630 26152 51686 26208
rect 51814 26424 51870 26480
rect 53010 27240 53066 27296
rect 53286 27512 53342 27568
rect 53194 27276 53196 27296
rect 53196 27276 53248 27296
rect 53248 27276 53250 27296
rect 53194 27240 53250 27276
rect 53102 27104 53158 27160
rect 54022 27240 54078 27296
rect 51998 2080 52054 2136
rect 55310 27276 55312 27296
rect 55312 27276 55364 27296
rect 55364 27276 55366 27296
rect 55310 27240 55366 27276
rect 57058 27784 57114 27840
rect 56414 27276 56416 27296
rect 56416 27276 56468 27296
rect 56468 27276 56470 27296
rect 56414 27240 56470 27276
rect 57702 27240 57758 27296
rect 57242 26696 57298 26752
rect 53838 2080 53894 2136
rect 55310 2080 55366 2136
rect 55218 1964 55274 2000
rect 55218 1944 55220 1964
rect 55220 1944 55272 1964
rect 55272 1944 55274 1964
rect 55586 2896 55642 2952
rect 55494 2624 55550 2680
rect 59542 27104 59598 27160
rect 59174 26560 59230 26616
rect 58438 26288 58494 26344
rect 57242 3168 57298 3224
rect 57978 3712 58034 3768
rect 58070 3596 58126 3632
rect 58070 3576 58072 3596
rect 58072 3576 58124 3596
rect 58124 3576 58126 3596
rect 58530 3576 58586 3632
rect 58070 3188 58126 3224
rect 58070 3168 58072 3188
rect 58072 3168 58124 3188
rect 58124 3168 58126 3188
rect 57702 3052 57758 3088
rect 57702 3032 57704 3052
rect 57704 3032 57756 3052
rect 57756 3032 57758 3052
rect 57794 2896 57850 2952
rect 57978 2796 57980 2816
rect 57980 2796 58032 2816
rect 58032 2796 58034 2816
rect 57978 2760 58034 2796
rect 58714 2896 58770 2952
rect 58806 2796 58808 2816
rect 58808 2796 58860 2816
rect 58860 2796 58862 2816
rect 58806 2760 58862 2796
rect 58162 1828 58218 1864
rect 58162 1808 58164 1828
rect 58164 1808 58216 1828
rect 58216 1808 58218 1828
rect 58070 1692 58126 1728
rect 58070 1672 58072 1692
rect 58072 1672 58124 1692
rect 58124 1672 58126 1692
rect 59852 27226 59908 27228
rect 59932 27226 59988 27228
rect 60012 27226 60068 27228
rect 60092 27226 60148 27228
rect 59852 27174 59898 27226
rect 59898 27174 59908 27226
rect 59932 27174 59962 27226
rect 59962 27174 59974 27226
rect 59974 27174 59988 27226
rect 60012 27174 60026 27226
rect 60026 27174 60038 27226
rect 60038 27174 60068 27226
rect 60092 27174 60102 27226
rect 60102 27174 60148 27226
rect 59852 27172 59908 27174
rect 59932 27172 59988 27174
rect 60012 27172 60068 27174
rect 60092 27172 60148 27174
rect 60646 27648 60702 27704
rect 60830 27648 60886 27704
rect 59726 26560 59782 26616
rect 59852 26138 59908 26140
rect 59932 26138 59988 26140
rect 60012 26138 60068 26140
rect 60092 26138 60148 26140
rect 59852 26086 59898 26138
rect 59898 26086 59908 26138
rect 59932 26086 59962 26138
rect 59962 26086 59974 26138
rect 59974 26086 59988 26138
rect 60012 26086 60026 26138
rect 60026 26086 60038 26138
rect 60038 26086 60068 26138
rect 60092 26086 60102 26138
rect 60102 26086 60148 26138
rect 59852 26084 59908 26086
rect 59932 26084 59988 26086
rect 60012 26084 60068 26086
rect 60092 26084 60148 26086
rect 60922 27532 60978 27568
rect 60922 27512 60924 27532
rect 60924 27512 60976 27532
rect 60976 27512 60978 27532
rect 60922 27240 60978 27296
rect 60738 27104 60794 27160
rect 60370 26696 60426 26752
rect 60554 26696 60610 26752
rect 60554 26424 60610 26480
rect 60646 26288 60702 26344
rect 60922 26560 60978 26616
rect 59634 25880 59690 25936
rect 61750 27512 61806 27568
rect 62302 27104 62358 27160
rect 61198 26424 61254 26480
rect 61750 26444 61806 26480
rect 61750 26424 61752 26444
rect 61752 26424 61804 26444
rect 61804 26424 61806 26444
rect 62302 26696 62358 26752
rect 62486 26696 62542 26752
rect 62210 26288 62266 26344
rect 59852 25050 59908 25052
rect 59932 25050 59988 25052
rect 60012 25050 60068 25052
rect 60092 25050 60148 25052
rect 59852 24998 59898 25050
rect 59898 24998 59908 25050
rect 59932 24998 59962 25050
rect 59962 24998 59974 25050
rect 59974 24998 59988 25050
rect 60012 24998 60026 25050
rect 60026 24998 60038 25050
rect 60038 24998 60068 25050
rect 60092 24998 60102 25050
rect 60102 24998 60148 25050
rect 59852 24996 59908 24998
rect 59932 24996 59988 24998
rect 60012 24996 60068 24998
rect 60092 24996 60148 24998
rect 59852 23962 59908 23964
rect 59932 23962 59988 23964
rect 60012 23962 60068 23964
rect 60092 23962 60148 23964
rect 59852 23910 59898 23962
rect 59898 23910 59908 23962
rect 59932 23910 59962 23962
rect 59962 23910 59974 23962
rect 59974 23910 59988 23962
rect 60012 23910 60026 23962
rect 60026 23910 60038 23962
rect 60038 23910 60068 23962
rect 60092 23910 60102 23962
rect 60102 23910 60148 23962
rect 59852 23908 59908 23910
rect 59932 23908 59988 23910
rect 60012 23908 60068 23910
rect 60092 23908 60148 23910
rect 59852 22874 59908 22876
rect 59932 22874 59988 22876
rect 60012 22874 60068 22876
rect 60092 22874 60148 22876
rect 59852 22822 59898 22874
rect 59898 22822 59908 22874
rect 59932 22822 59962 22874
rect 59962 22822 59974 22874
rect 59974 22822 59988 22874
rect 60012 22822 60026 22874
rect 60026 22822 60038 22874
rect 60038 22822 60068 22874
rect 60092 22822 60102 22874
rect 60102 22822 60148 22874
rect 59852 22820 59908 22822
rect 59932 22820 59988 22822
rect 60012 22820 60068 22822
rect 60092 22820 60148 22822
rect 59852 21786 59908 21788
rect 59932 21786 59988 21788
rect 60012 21786 60068 21788
rect 60092 21786 60148 21788
rect 59852 21734 59898 21786
rect 59898 21734 59908 21786
rect 59932 21734 59962 21786
rect 59962 21734 59974 21786
rect 59974 21734 59988 21786
rect 60012 21734 60026 21786
rect 60026 21734 60038 21786
rect 60038 21734 60068 21786
rect 60092 21734 60102 21786
rect 60102 21734 60148 21786
rect 59852 21732 59908 21734
rect 59932 21732 59988 21734
rect 60012 21732 60068 21734
rect 60092 21732 60148 21734
rect 59852 20698 59908 20700
rect 59932 20698 59988 20700
rect 60012 20698 60068 20700
rect 60092 20698 60148 20700
rect 59852 20646 59898 20698
rect 59898 20646 59908 20698
rect 59932 20646 59962 20698
rect 59962 20646 59974 20698
rect 59974 20646 59988 20698
rect 60012 20646 60026 20698
rect 60026 20646 60038 20698
rect 60038 20646 60068 20698
rect 60092 20646 60102 20698
rect 60102 20646 60148 20698
rect 59852 20644 59908 20646
rect 59932 20644 59988 20646
rect 60012 20644 60068 20646
rect 60092 20644 60148 20646
rect 59852 19610 59908 19612
rect 59932 19610 59988 19612
rect 60012 19610 60068 19612
rect 60092 19610 60148 19612
rect 59852 19558 59898 19610
rect 59898 19558 59908 19610
rect 59932 19558 59962 19610
rect 59962 19558 59974 19610
rect 59974 19558 59988 19610
rect 60012 19558 60026 19610
rect 60026 19558 60038 19610
rect 60038 19558 60068 19610
rect 60092 19558 60102 19610
rect 60102 19558 60148 19610
rect 59852 19556 59908 19558
rect 59932 19556 59988 19558
rect 60012 19556 60068 19558
rect 60092 19556 60148 19558
rect 59852 18522 59908 18524
rect 59932 18522 59988 18524
rect 60012 18522 60068 18524
rect 60092 18522 60148 18524
rect 59852 18470 59898 18522
rect 59898 18470 59908 18522
rect 59932 18470 59962 18522
rect 59962 18470 59974 18522
rect 59974 18470 59988 18522
rect 60012 18470 60026 18522
rect 60026 18470 60038 18522
rect 60038 18470 60068 18522
rect 60092 18470 60102 18522
rect 60102 18470 60148 18522
rect 59852 18468 59908 18470
rect 59932 18468 59988 18470
rect 60012 18468 60068 18470
rect 60092 18468 60148 18470
rect 59852 17434 59908 17436
rect 59932 17434 59988 17436
rect 60012 17434 60068 17436
rect 60092 17434 60148 17436
rect 59852 17382 59898 17434
rect 59898 17382 59908 17434
rect 59932 17382 59962 17434
rect 59962 17382 59974 17434
rect 59974 17382 59988 17434
rect 60012 17382 60026 17434
rect 60026 17382 60038 17434
rect 60038 17382 60068 17434
rect 60092 17382 60102 17434
rect 60102 17382 60148 17434
rect 59852 17380 59908 17382
rect 59932 17380 59988 17382
rect 60012 17380 60068 17382
rect 60092 17380 60148 17382
rect 59634 3732 59690 3768
rect 59634 3712 59636 3732
rect 59636 3712 59688 3732
rect 59688 3712 59690 3732
rect 59852 16346 59908 16348
rect 59932 16346 59988 16348
rect 60012 16346 60068 16348
rect 60092 16346 60148 16348
rect 59852 16294 59898 16346
rect 59898 16294 59908 16346
rect 59932 16294 59962 16346
rect 59962 16294 59974 16346
rect 59974 16294 59988 16346
rect 60012 16294 60026 16346
rect 60026 16294 60038 16346
rect 60038 16294 60068 16346
rect 60092 16294 60102 16346
rect 60102 16294 60148 16346
rect 59852 16292 59908 16294
rect 59932 16292 59988 16294
rect 60012 16292 60068 16294
rect 60092 16292 60148 16294
rect 59852 15258 59908 15260
rect 59932 15258 59988 15260
rect 60012 15258 60068 15260
rect 60092 15258 60148 15260
rect 59852 15206 59898 15258
rect 59898 15206 59908 15258
rect 59932 15206 59962 15258
rect 59962 15206 59974 15258
rect 59974 15206 59988 15258
rect 60012 15206 60026 15258
rect 60026 15206 60038 15258
rect 60038 15206 60068 15258
rect 60092 15206 60102 15258
rect 60102 15206 60148 15258
rect 59852 15204 59908 15206
rect 59932 15204 59988 15206
rect 60012 15204 60068 15206
rect 60092 15204 60148 15206
rect 59852 14170 59908 14172
rect 59932 14170 59988 14172
rect 60012 14170 60068 14172
rect 60092 14170 60148 14172
rect 59852 14118 59898 14170
rect 59898 14118 59908 14170
rect 59932 14118 59962 14170
rect 59962 14118 59974 14170
rect 59974 14118 59988 14170
rect 60012 14118 60026 14170
rect 60026 14118 60038 14170
rect 60038 14118 60068 14170
rect 60092 14118 60102 14170
rect 60102 14118 60148 14170
rect 59852 14116 59908 14118
rect 59932 14116 59988 14118
rect 60012 14116 60068 14118
rect 60092 14116 60148 14118
rect 59852 13082 59908 13084
rect 59932 13082 59988 13084
rect 60012 13082 60068 13084
rect 60092 13082 60148 13084
rect 59852 13030 59898 13082
rect 59898 13030 59908 13082
rect 59932 13030 59962 13082
rect 59962 13030 59974 13082
rect 59974 13030 59988 13082
rect 60012 13030 60026 13082
rect 60026 13030 60038 13082
rect 60038 13030 60068 13082
rect 60092 13030 60102 13082
rect 60102 13030 60148 13082
rect 59852 13028 59908 13030
rect 59932 13028 59988 13030
rect 60012 13028 60068 13030
rect 60092 13028 60148 13030
rect 59852 11994 59908 11996
rect 59932 11994 59988 11996
rect 60012 11994 60068 11996
rect 60092 11994 60148 11996
rect 59852 11942 59898 11994
rect 59898 11942 59908 11994
rect 59932 11942 59962 11994
rect 59962 11942 59974 11994
rect 59974 11942 59988 11994
rect 60012 11942 60026 11994
rect 60026 11942 60038 11994
rect 60038 11942 60068 11994
rect 60092 11942 60102 11994
rect 60102 11942 60148 11994
rect 59852 11940 59908 11942
rect 59932 11940 59988 11942
rect 60012 11940 60068 11942
rect 60092 11940 60148 11942
rect 59852 10906 59908 10908
rect 59932 10906 59988 10908
rect 60012 10906 60068 10908
rect 60092 10906 60148 10908
rect 59852 10854 59898 10906
rect 59898 10854 59908 10906
rect 59932 10854 59962 10906
rect 59962 10854 59974 10906
rect 59974 10854 59988 10906
rect 60012 10854 60026 10906
rect 60026 10854 60038 10906
rect 60038 10854 60068 10906
rect 60092 10854 60102 10906
rect 60102 10854 60148 10906
rect 59852 10852 59908 10854
rect 59932 10852 59988 10854
rect 60012 10852 60068 10854
rect 60092 10852 60148 10854
rect 59852 9818 59908 9820
rect 59932 9818 59988 9820
rect 60012 9818 60068 9820
rect 60092 9818 60148 9820
rect 59852 9766 59898 9818
rect 59898 9766 59908 9818
rect 59932 9766 59962 9818
rect 59962 9766 59974 9818
rect 59974 9766 59988 9818
rect 60012 9766 60026 9818
rect 60026 9766 60038 9818
rect 60038 9766 60068 9818
rect 60092 9766 60102 9818
rect 60102 9766 60148 9818
rect 59852 9764 59908 9766
rect 59932 9764 59988 9766
rect 60012 9764 60068 9766
rect 60092 9764 60148 9766
rect 59852 8730 59908 8732
rect 59932 8730 59988 8732
rect 60012 8730 60068 8732
rect 60092 8730 60148 8732
rect 59852 8678 59898 8730
rect 59898 8678 59908 8730
rect 59932 8678 59962 8730
rect 59962 8678 59974 8730
rect 59974 8678 59988 8730
rect 60012 8678 60026 8730
rect 60026 8678 60038 8730
rect 60038 8678 60068 8730
rect 60092 8678 60102 8730
rect 60102 8678 60148 8730
rect 59852 8676 59908 8678
rect 59932 8676 59988 8678
rect 60012 8676 60068 8678
rect 60092 8676 60148 8678
rect 59852 7642 59908 7644
rect 59932 7642 59988 7644
rect 60012 7642 60068 7644
rect 60092 7642 60148 7644
rect 59852 7590 59898 7642
rect 59898 7590 59908 7642
rect 59932 7590 59962 7642
rect 59962 7590 59974 7642
rect 59974 7590 59988 7642
rect 60012 7590 60026 7642
rect 60026 7590 60038 7642
rect 60038 7590 60068 7642
rect 60092 7590 60102 7642
rect 60102 7590 60148 7642
rect 59852 7588 59908 7590
rect 59932 7588 59988 7590
rect 60012 7588 60068 7590
rect 60092 7588 60148 7590
rect 59852 6554 59908 6556
rect 59932 6554 59988 6556
rect 60012 6554 60068 6556
rect 60092 6554 60148 6556
rect 59852 6502 59898 6554
rect 59898 6502 59908 6554
rect 59932 6502 59962 6554
rect 59962 6502 59974 6554
rect 59974 6502 59988 6554
rect 60012 6502 60026 6554
rect 60026 6502 60038 6554
rect 60038 6502 60068 6554
rect 60092 6502 60102 6554
rect 60102 6502 60148 6554
rect 59852 6500 59908 6502
rect 59932 6500 59988 6502
rect 60012 6500 60068 6502
rect 60092 6500 60148 6502
rect 59852 5466 59908 5468
rect 59932 5466 59988 5468
rect 60012 5466 60068 5468
rect 60092 5466 60148 5468
rect 59852 5414 59898 5466
rect 59898 5414 59908 5466
rect 59932 5414 59962 5466
rect 59962 5414 59974 5466
rect 59974 5414 59988 5466
rect 60012 5414 60026 5466
rect 60026 5414 60038 5466
rect 60038 5414 60068 5466
rect 60092 5414 60102 5466
rect 60102 5414 60148 5466
rect 59852 5412 59908 5414
rect 59932 5412 59988 5414
rect 60012 5412 60068 5414
rect 60092 5412 60148 5414
rect 59852 4378 59908 4380
rect 59932 4378 59988 4380
rect 60012 4378 60068 4380
rect 60092 4378 60148 4380
rect 59852 4326 59898 4378
rect 59898 4326 59908 4378
rect 59932 4326 59962 4378
rect 59962 4326 59974 4378
rect 59974 4326 59988 4378
rect 60012 4326 60026 4378
rect 60026 4326 60038 4378
rect 60038 4326 60068 4378
rect 60092 4326 60102 4378
rect 60102 4326 60148 4378
rect 59852 4324 59908 4326
rect 59932 4324 59988 4326
rect 60012 4324 60068 4326
rect 60092 4324 60148 4326
rect 59852 3290 59908 3292
rect 59932 3290 59988 3292
rect 60012 3290 60068 3292
rect 60092 3290 60148 3292
rect 59852 3238 59898 3290
rect 59898 3238 59908 3290
rect 59932 3238 59962 3290
rect 59962 3238 59974 3290
rect 59974 3238 59988 3290
rect 60012 3238 60026 3290
rect 60026 3238 60038 3290
rect 60038 3238 60068 3290
rect 60092 3238 60102 3290
rect 60102 3238 60148 3290
rect 59852 3236 59908 3238
rect 59932 3236 59988 3238
rect 60012 3236 60068 3238
rect 60092 3236 60148 3238
rect 59852 2202 59908 2204
rect 59932 2202 59988 2204
rect 60012 2202 60068 2204
rect 60092 2202 60148 2204
rect 59852 2150 59898 2202
rect 59898 2150 59908 2202
rect 59932 2150 59962 2202
rect 59962 2150 59974 2202
rect 59974 2150 59988 2202
rect 60012 2150 60026 2202
rect 60026 2150 60038 2202
rect 60038 2150 60068 2202
rect 60092 2150 60102 2202
rect 60102 2150 60148 2202
rect 59852 2148 59908 2150
rect 59932 2148 59988 2150
rect 60012 2148 60068 2150
rect 60092 2148 60148 2150
rect 60922 2760 60978 2816
rect 60646 2100 60702 2136
rect 60646 2080 60648 2100
rect 60648 2080 60700 2100
rect 60700 2080 60702 2100
rect 61014 2252 61016 2272
rect 61016 2252 61068 2272
rect 61068 2252 61070 2272
rect 61014 2216 61070 2252
rect 61014 1980 61016 2000
rect 61016 1980 61068 2000
rect 61068 1980 61070 2000
rect 61014 1944 61070 1980
rect 60830 1672 60886 1728
rect 61290 1672 61346 1728
rect 63222 26152 63278 26208
rect 65062 26424 65118 26480
rect 62578 2624 62634 2680
rect 62762 2644 62818 2680
rect 62762 2624 62764 2644
rect 62764 2624 62816 2644
rect 62816 2624 62818 2644
rect 64050 2896 64106 2952
rect 68374 27240 68430 27296
rect 64142 1672 64198 1728
rect 66166 3032 66222 3088
rect 69018 25880 69074 25936
rect 68650 14884 68706 14920
rect 68650 14864 68652 14884
rect 68652 14864 68704 14884
rect 68704 14864 68706 14884
rect 69938 27784 69994 27840
rect 69570 26732 69572 26752
rect 69572 26732 69624 26752
rect 69624 26732 69626 26752
rect 69570 26696 69626 26732
rect 69846 26696 69902 26752
rect 70490 26696 70546 26752
rect 70490 26152 70546 26208
rect 67270 2624 67326 2680
rect 67454 2080 67510 2136
rect 67362 1808 67418 1864
rect 66902 1692 66958 1728
rect 66902 1672 66904 1692
rect 66904 1672 66956 1692
rect 66956 1672 66958 1692
rect 70214 14884 70270 14920
rect 70214 14864 70216 14884
rect 70216 14864 70268 14884
rect 70268 14864 70270 14884
rect 69938 2216 69994 2272
rect 70306 3068 70308 3088
rect 70308 3068 70360 3088
rect 70360 3068 70362 3088
rect 70306 3032 70362 3068
rect 70674 2216 70730 2272
rect 71870 26188 71872 26208
rect 71872 26188 71924 26208
rect 71924 26188 71926 26208
rect 71870 26152 71926 26188
rect 72422 27240 72478 27296
rect 72238 26560 72294 26616
rect 72514 25880 72570 25936
rect 74906 27920 74962 27976
rect 73802 27784 73858 27840
rect 73066 26732 73068 26752
rect 73068 26732 73120 26752
rect 73120 26732 73122 26752
rect 73066 26696 73122 26732
rect 70950 1844 70952 1864
rect 70952 1844 71004 1864
rect 71004 1844 71006 1864
rect 70950 1808 71006 1844
rect 72330 1944 72386 2000
rect 74576 27770 74632 27772
rect 74656 27770 74712 27772
rect 74736 27770 74792 27772
rect 74816 27770 74872 27772
rect 74576 27718 74622 27770
rect 74622 27718 74632 27770
rect 74656 27718 74686 27770
rect 74686 27718 74698 27770
rect 74698 27718 74712 27770
rect 74736 27718 74750 27770
rect 74750 27718 74762 27770
rect 74762 27718 74792 27770
rect 74816 27718 74826 27770
rect 74826 27718 74872 27770
rect 74576 27716 74632 27718
rect 74656 27716 74712 27718
rect 74736 27716 74792 27718
rect 74816 27716 74872 27718
rect 74262 27648 74318 27704
rect 74814 27104 74870 27160
rect 74576 26682 74632 26684
rect 74656 26682 74712 26684
rect 74736 26682 74792 26684
rect 74816 26682 74872 26684
rect 74576 26630 74622 26682
rect 74622 26630 74632 26682
rect 74656 26630 74686 26682
rect 74686 26630 74698 26682
rect 74698 26630 74712 26682
rect 74736 26630 74750 26682
rect 74750 26630 74762 26682
rect 74762 26630 74792 26682
rect 74816 26630 74826 26682
rect 74826 26630 74872 26682
rect 74576 26628 74632 26630
rect 74656 26628 74712 26630
rect 74736 26628 74792 26630
rect 74816 26628 74872 26630
rect 75182 27648 75238 27704
rect 75550 26832 75606 26888
rect 76562 27104 76618 27160
rect 74576 25594 74632 25596
rect 74656 25594 74712 25596
rect 74736 25594 74792 25596
rect 74816 25594 74872 25596
rect 74576 25542 74622 25594
rect 74622 25542 74632 25594
rect 74656 25542 74686 25594
rect 74686 25542 74698 25594
rect 74698 25542 74712 25594
rect 74736 25542 74750 25594
rect 74750 25542 74762 25594
rect 74762 25542 74792 25594
rect 74816 25542 74826 25594
rect 74826 25542 74872 25594
rect 74576 25540 74632 25542
rect 74656 25540 74712 25542
rect 74736 25540 74792 25542
rect 74816 25540 74872 25542
rect 74576 24506 74632 24508
rect 74656 24506 74712 24508
rect 74736 24506 74792 24508
rect 74816 24506 74872 24508
rect 74576 24454 74622 24506
rect 74622 24454 74632 24506
rect 74656 24454 74686 24506
rect 74686 24454 74698 24506
rect 74698 24454 74712 24506
rect 74736 24454 74750 24506
rect 74750 24454 74762 24506
rect 74762 24454 74792 24506
rect 74816 24454 74826 24506
rect 74826 24454 74872 24506
rect 74576 24452 74632 24454
rect 74656 24452 74712 24454
rect 74736 24452 74792 24454
rect 74816 24452 74872 24454
rect 74576 23418 74632 23420
rect 74656 23418 74712 23420
rect 74736 23418 74792 23420
rect 74816 23418 74872 23420
rect 74576 23366 74622 23418
rect 74622 23366 74632 23418
rect 74656 23366 74686 23418
rect 74686 23366 74698 23418
rect 74698 23366 74712 23418
rect 74736 23366 74750 23418
rect 74750 23366 74762 23418
rect 74762 23366 74792 23418
rect 74816 23366 74826 23418
rect 74826 23366 74872 23418
rect 74576 23364 74632 23366
rect 74656 23364 74712 23366
rect 74736 23364 74792 23366
rect 74816 23364 74872 23366
rect 74576 22330 74632 22332
rect 74656 22330 74712 22332
rect 74736 22330 74792 22332
rect 74816 22330 74872 22332
rect 74576 22278 74622 22330
rect 74622 22278 74632 22330
rect 74656 22278 74686 22330
rect 74686 22278 74698 22330
rect 74698 22278 74712 22330
rect 74736 22278 74750 22330
rect 74750 22278 74762 22330
rect 74762 22278 74792 22330
rect 74816 22278 74826 22330
rect 74826 22278 74872 22330
rect 74576 22276 74632 22278
rect 74656 22276 74712 22278
rect 74736 22276 74792 22278
rect 74816 22276 74872 22278
rect 74576 21242 74632 21244
rect 74656 21242 74712 21244
rect 74736 21242 74792 21244
rect 74816 21242 74872 21244
rect 74576 21190 74622 21242
rect 74622 21190 74632 21242
rect 74656 21190 74686 21242
rect 74686 21190 74698 21242
rect 74698 21190 74712 21242
rect 74736 21190 74750 21242
rect 74750 21190 74762 21242
rect 74762 21190 74792 21242
rect 74816 21190 74826 21242
rect 74826 21190 74872 21242
rect 74576 21188 74632 21190
rect 74656 21188 74712 21190
rect 74736 21188 74792 21190
rect 74816 21188 74872 21190
rect 74576 20154 74632 20156
rect 74656 20154 74712 20156
rect 74736 20154 74792 20156
rect 74816 20154 74872 20156
rect 74576 20102 74622 20154
rect 74622 20102 74632 20154
rect 74656 20102 74686 20154
rect 74686 20102 74698 20154
rect 74698 20102 74712 20154
rect 74736 20102 74750 20154
rect 74750 20102 74762 20154
rect 74762 20102 74792 20154
rect 74816 20102 74826 20154
rect 74826 20102 74872 20154
rect 74576 20100 74632 20102
rect 74656 20100 74712 20102
rect 74736 20100 74792 20102
rect 74816 20100 74872 20102
rect 74576 19066 74632 19068
rect 74656 19066 74712 19068
rect 74736 19066 74792 19068
rect 74816 19066 74872 19068
rect 74576 19014 74622 19066
rect 74622 19014 74632 19066
rect 74656 19014 74686 19066
rect 74686 19014 74698 19066
rect 74698 19014 74712 19066
rect 74736 19014 74750 19066
rect 74750 19014 74762 19066
rect 74762 19014 74792 19066
rect 74816 19014 74826 19066
rect 74826 19014 74872 19066
rect 74576 19012 74632 19014
rect 74656 19012 74712 19014
rect 74736 19012 74792 19014
rect 74816 19012 74872 19014
rect 74576 17978 74632 17980
rect 74656 17978 74712 17980
rect 74736 17978 74792 17980
rect 74816 17978 74872 17980
rect 74576 17926 74622 17978
rect 74622 17926 74632 17978
rect 74656 17926 74686 17978
rect 74686 17926 74698 17978
rect 74698 17926 74712 17978
rect 74736 17926 74750 17978
rect 74750 17926 74762 17978
rect 74762 17926 74792 17978
rect 74816 17926 74826 17978
rect 74826 17926 74872 17978
rect 74576 17924 74632 17926
rect 74656 17924 74712 17926
rect 74736 17924 74792 17926
rect 74816 17924 74872 17926
rect 74576 16890 74632 16892
rect 74656 16890 74712 16892
rect 74736 16890 74792 16892
rect 74816 16890 74872 16892
rect 74576 16838 74622 16890
rect 74622 16838 74632 16890
rect 74656 16838 74686 16890
rect 74686 16838 74698 16890
rect 74698 16838 74712 16890
rect 74736 16838 74750 16890
rect 74750 16838 74762 16890
rect 74762 16838 74792 16890
rect 74816 16838 74826 16890
rect 74826 16838 74872 16890
rect 74576 16836 74632 16838
rect 74656 16836 74712 16838
rect 74736 16836 74792 16838
rect 74816 16836 74872 16838
rect 74576 15802 74632 15804
rect 74656 15802 74712 15804
rect 74736 15802 74792 15804
rect 74816 15802 74872 15804
rect 74576 15750 74622 15802
rect 74622 15750 74632 15802
rect 74656 15750 74686 15802
rect 74686 15750 74698 15802
rect 74698 15750 74712 15802
rect 74736 15750 74750 15802
rect 74750 15750 74762 15802
rect 74762 15750 74792 15802
rect 74816 15750 74826 15802
rect 74826 15750 74872 15802
rect 74576 15748 74632 15750
rect 74656 15748 74712 15750
rect 74736 15748 74792 15750
rect 74816 15748 74872 15750
rect 74576 14714 74632 14716
rect 74656 14714 74712 14716
rect 74736 14714 74792 14716
rect 74816 14714 74872 14716
rect 74576 14662 74622 14714
rect 74622 14662 74632 14714
rect 74656 14662 74686 14714
rect 74686 14662 74698 14714
rect 74698 14662 74712 14714
rect 74736 14662 74750 14714
rect 74750 14662 74762 14714
rect 74762 14662 74792 14714
rect 74816 14662 74826 14714
rect 74826 14662 74872 14714
rect 74576 14660 74632 14662
rect 74656 14660 74712 14662
rect 74736 14660 74792 14662
rect 74816 14660 74872 14662
rect 74576 13626 74632 13628
rect 74656 13626 74712 13628
rect 74736 13626 74792 13628
rect 74816 13626 74872 13628
rect 74576 13574 74622 13626
rect 74622 13574 74632 13626
rect 74656 13574 74686 13626
rect 74686 13574 74698 13626
rect 74698 13574 74712 13626
rect 74736 13574 74750 13626
rect 74750 13574 74762 13626
rect 74762 13574 74792 13626
rect 74816 13574 74826 13626
rect 74826 13574 74872 13626
rect 74576 13572 74632 13574
rect 74656 13572 74712 13574
rect 74736 13572 74792 13574
rect 74816 13572 74872 13574
rect 74576 12538 74632 12540
rect 74656 12538 74712 12540
rect 74736 12538 74792 12540
rect 74816 12538 74872 12540
rect 74576 12486 74622 12538
rect 74622 12486 74632 12538
rect 74656 12486 74686 12538
rect 74686 12486 74698 12538
rect 74698 12486 74712 12538
rect 74736 12486 74750 12538
rect 74750 12486 74762 12538
rect 74762 12486 74792 12538
rect 74816 12486 74826 12538
rect 74826 12486 74872 12538
rect 74576 12484 74632 12486
rect 74656 12484 74712 12486
rect 74736 12484 74792 12486
rect 74816 12484 74872 12486
rect 74576 11450 74632 11452
rect 74656 11450 74712 11452
rect 74736 11450 74792 11452
rect 74816 11450 74872 11452
rect 74576 11398 74622 11450
rect 74622 11398 74632 11450
rect 74656 11398 74686 11450
rect 74686 11398 74698 11450
rect 74698 11398 74712 11450
rect 74736 11398 74750 11450
rect 74750 11398 74762 11450
rect 74762 11398 74792 11450
rect 74816 11398 74826 11450
rect 74826 11398 74872 11450
rect 74576 11396 74632 11398
rect 74656 11396 74712 11398
rect 74736 11396 74792 11398
rect 74816 11396 74872 11398
rect 74576 10362 74632 10364
rect 74656 10362 74712 10364
rect 74736 10362 74792 10364
rect 74816 10362 74872 10364
rect 74576 10310 74622 10362
rect 74622 10310 74632 10362
rect 74656 10310 74686 10362
rect 74686 10310 74698 10362
rect 74698 10310 74712 10362
rect 74736 10310 74750 10362
rect 74750 10310 74762 10362
rect 74762 10310 74792 10362
rect 74816 10310 74826 10362
rect 74826 10310 74872 10362
rect 74576 10308 74632 10310
rect 74656 10308 74712 10310
rect 74736 10308 74792 10310
rect 74816 10308 74872 10310
rect 74576 9274 74632 9276
rect 74656 9274 74712 9276
rect 74736 9274 74792 9276
rect 74816 9274 74872 9276
rect 74576 9222 74622 9274
rect 74622 9222 74632 9274
rect 74656 9222 74686 9274
rect 74686 9222 74698 9274
rect 74698 9222 74712 9274
rect 74736 9222 74750 9274
rect 74750 9222 74762 9274
rect 74762 9222 74792 9274
rect 74816 9222 74826 9274
rect 74826 9222 74872 9274
rect 74576 9220 74632 9222
rect 74656 9220 74712 9222
rect 74736 9220 74792 9222
rect 74816 9220 74872 9222
rect 74576 8186 74632 8188
rect 74656 8186 74712 8188
rect 74736 8186 74792 8188
rect 74816 8186 74872 8188
rect 74576 8134 74622 8186
rect 74622 8134 74632 8186
rect 74656 8134 74686 8186
rect 74686 8134 74698 8186
rect 74698 8134 74712 8186
rect 74736 8134 74750 8186
rect 74750 8134 74762 8186
rect 74762 8134 74792 8186
rect 74816 8134 74826 8186
rect 74826 8134 74872 8186
rect 74576 8132 74632 8134
rect 74656 8132 74712 8134
rect 74736 8132 74792 8134
rect 74816 8132 74872 8134
rect 74576 7098 74632 7100
rect 74656 7098 74712 7100
rect 74736 7098 74792 7100
rect 74816 7098 74872 7100
rect 74576 7046 74622 7098
rect 74622 7046 74632 7098
rect 74656 7046 74686 7098
rect 74686 7046 74698 7098
rect 74698 7046 74712 7098
rect 74736 7046 74750 7098
rect 74750 7046 74762 7098
rect 74762 7046 74792 7098
rect 74816 7046 74826 7098
rect 74826 7046 74872 7098
rect 74576 7044 74632 7046
rect 74656 7044 74712 7046
rect 74736 7044 74792 7046
rect 74816 7044 74872 7046
rect 74576 6010 74632 6012
rect 74656 6010 74712 6012
rect 74736 6010 74792 6012
rect 74816 6010 74872 6012
rect 74576 5958 74622 6010
rect 74622 5958 74632 6010
rect 74656 5958 74686 6010
rect 74686 5958 74698 6010
rect 74698 5958 74712 6010
rect 74736 5958 74750 6010
rect 74750 5958 74762 6010
rect 74762 5958 74792 6010
rect 74816 5958 74826 6010
rect 74826 5958 74872 6010
rect 74576 5956 74632 5958
rect 74656 5956 74712 5958
rect 74736 5956 74792 5958
rect 74816 5956 74872 5958
rect 74576 4922 74632 4924
rect 74656 4922 74712 4924
rect 74736 4922 74792 4924
rect 74816 4922 74872 4924
rect 74576 4870 74622 4922
rect 74622 4870 74632 4922
rect 74656 4870 74686 4922
rect 74686 4870 74698 4922
rect 74698 4870 74712 4922
rect 74736 4870 74750 4922
rect 74750 4870 74762 4922
rect 74762 4870 74792 4922
rect 74816 4870 74826 4922
rect 74826 4870 74872 4922
rect 74576 4868 74632 4870
rect 74656 4868 74712 4870
rect 74736 4868 74792 4870
rect 74816 4868 74872 4870
rect 72882 1672 72938 1728
rect 73434 2796 73436 2816
rect 73436 2796 73488 2816
rect 73488 2796 73490 2816
rect 73434 2760 73490 2796
rect 74576 3834 74632 3836
rect 74656 3834 74712 3836
rect 74736 3834 74792 3836
rect 74816 3834 74872 3836
rect 74576 3782 74622 3834
rect 74622 3782 74632 3834
rect 74656 3782 74686 3834
rect 74686 3782 74698 3834
rect 74698 3782 74712 3834
rect 74736 3782 74750 3834
rect 74750 3782 74762 3834
rect 74762 3782 74792 3834
rect 74816 3782 74826 3834
rect 74826 3782 74872 3834
rect 74576 3780 74632 3782
rect 74656 3780 74712 3782
rect 74736 3780 74792 3782
rect 74816 3780 74872 3782
rect 74576 2746 74632 2748
rect 74656 2746 74712 2748
rect 74736 2746 74792 2748
rect 74816 2746 74872 2748
rect 74576 2694 74622 2746
rect 74622 2694 74632 2746
rect 74656 2694 74686 2746
rect 74686 2694 74698 2746
rect 74698 2694 74712 2746
rect 74736 2694 74750 2746
rect 74750 2694 74762 2746
rect 74762 2694 74792 2746
rect 74816 2694 74826 2746
rect 74826 2694 74872 2746
rect 74576 2692 74632 2694
rect 74656 2692 74712 2694
rect 74736 2692 74792 2694
rect 74816 2692 74872 2694
rect 74630 2488 74686 2544
rect 78586 27276 78588 27296
rect 78588 27276 78640 27296
rect 78640 27276 78642 27296
rect 78586 27240 78642 27276
rect 78770 26560 78826 26616
rect 79046 27376 79102 27432
rect 77114 3032 77170 3088
rect 79414 27648 79470 27704
rect 79322 27104 79378 27160
rect 80242 27240 80298 27296
rect 80334 27104 80390 27160
rect 80058 26832 80114 26888
rect 80242 26832 80298 26888
rect 79690 26424 79746 26480
rect 80242 26288 80298 26344
rect 81162 26696 81218 26752
rect 81898 26560 81954 26616
rect 81438 26424 81494 26480
rect 80426 26288 80482 26344
rect 77206 2760 77262 2816
rect 75550 1844 75552 1864
rect 75552 1844 75604 1864
rect 75604 1844 75606 1864
rect 75550 1808 75606 1844
rect 78034 2760 78090 2816
rect 79782 26152 79838 26208
rect 85210 27920 85266 27976
rect 84474 27276 84476 27296
rect 84476 27276 84528 27296
rect 84528 27276 84530 27296
rect 84474 27240 84530 27276
rect 77390 1944 77446 2000
rect 77850 1692 77906 1728
rect 77850 1672 77852 1692
rect 77852 1672 77904 1692
rect 77904 1672 77906 1692
rect 79598 2216 79654 2272
rect 80150 2216 80206 2272
rect 80058 1420 80114 1456
rect 80058 1400 80060 1420
rect 80060 1400 80112 1420
rect 80112 1400 80114 1420
rect 85210 27240 85266 27296
rect 89074 27376 89130 27432
rect 87326 27104 87382 27160
rect 89300 27226 89356 27228
rect 89380 27226 89436 27228
rect 89460 27226 89516 27228
rect 89540 27226 89596 27228
rect 89300 27174 89346 27226
rect 89346 27174 89356 27226
rect 89380 27174 89410 27226
rect 89410 27174 89422 27226
rect 89422 27174 89436 27226
rect 89460 27174 89474 27226
rect 89474 27174 89486 27226
rect 89486 27174 89516 27226
rect 89540 27174 89550 27226
rect 89550 27174 89596 27226
rect 89300 27172 89356 27174
rect 89380 27172 89436 27174
rect 89460 27172 89516 27174
rect 89540 27172 89596 27174
rect 89074 26424 89130 26480
rect 90362 27104 90418 27160
rect 89300 26138 89356 26140
rect 89380 26138 89436 26140
rect 89460 26138 89516 26140
rect 89540 26138 89596 26140
rect 89300 26086 89346 26138
rect 89346 26086 89356 26138
rect 89380 26086 89410 26138
rect 89410 26086 89422 26138
rect 89422 26086 89436 26138
rect 89460 26086 89474 26138
rect 89474 26086 89486 26138
rect 89486 26086 89516 26138
rect 89540 26086 89550 26138
rect 89550 26086 89596 26138
rect 89300 26084 89356 26086
rect 89380 26084 89436 26086
rect 89460 26084 89516 26086
rect 89540 26084 89596 26086
rect 89300 25050 89356 25052
rect 89380 25050 89436 25052
rect 89460 25050 89516 25052
rect 89540 25050 89596 25052
rect 89300 24998 89346 25050
rect 89346 24998 89356 25050
rect 89380 24998 89410 25050
rect 89410 24998 89422 25050
rect 89422 24998 89436 25050
rect 89460 24998 89474 25050
rect 89474 24998 89486 25050
rect 89486 24998 89516 25050
rect 89540 24998 89550 25050
rect 89550 24998 89596 25050
rect 89300 24996 89356 24998
rect 89380 24996 89436 24998
rect 89460 24996 89516 24998
rect 89540 24996 89596 24998
rect 89300 23962 89356 23964
rect 89380 23962 89436 23964
rect 89460 23962 89516 23964
rect 89540 23962 89596 23964
rect 89300 23910 89346 23962
rect 89346 23910 89356 23962
rect 89380 23910 89410 23962
rect 89410 23910 89422 23962
rect 89422 23910 89436 23962
rect 89460 23910 89474 23962
rect 89474 23910 89486 23962
rect 89486 23910 89516 23962
rect 89540 23910 89550 23962
rect 89550 23910 89596 23962
rect 89300 23908 89356 23910
rect 89380 23908 89436 23910
rect 89460 23908 89516 23910
rect 89540 23908 89596 23910
rect 89300 22874 89356 22876
rect 89380 22874 89436 22876
rect 89460 22874 89516 22876
rect 89540 22874 89596 22876
rect 89300 22822 89346 22874
rect 89346 22822 89356 22874
rect 89380 22822 89410 22874
rect 89410 22822 89422 22874
rect 89422 22822 89436 22874
rect 89460 22822 89474 22874
rect 89474 22822 89486 22874
rect 89486 22822 89516 22874
rect 89540 22822 89550 22874
rect 89550 22822 89596 22874
rect 89300 22820 89356 22822
rect 89380 22820 89436 22822
rect 89460 22820 89516 22822
rect 89540 22820 89596 22822
rect 89300 21786 89356 21788
rect 89380 21786 89436 21788
rect 89460 21786 89516 21788
rect 89540 21786 89596 21788
rect 89300 21734 89346 21786
rect 89346 21734 89356 21786
rect 89380 21734 89410 21786
rect 89410 21734 89422 21786
rect 89422 21734 89436 21786
rect 89460 21734 89474 21786
rect 89474 21734 89486 21786
rect 89486 21734 89516 21786
rect 89540 21734 89550 21786
rect 89550 21734 89596 21786
rect 89300 21732 89356 21734
rect 89380 21732 89436 21734
rect 89460 21732 89516 21734
rect 89540 21732 89596 21734
rect 89300 20698 89356 20700
rect 89380 20698 89436 20700
rect 89460 20698 89516 20700
rect 89540 20698 89596 20700
rect 89300 20646 89346 20698
rect 89346 20646 89356 20698
rect 89380 20646 89410 20698
rect 89410 20646 89422 20698
rect 89422 20646 89436 20698
rect 89460 20646 89474 20698
rect 89474 20646 89486 20698
rect 89486 20646 89516 20698
rect 89540 20646 89550 20698
rect 89550 20646 89596 20698
rect 89300 20644 89356 20646
rect 89380 20644 89436 20646
rect 89460 20644 89516 20646
rect 89540 20644 89596 20646
rect 89300 19610 89356 19612
rect 89380 19610 89436 19612
rect 89460 19610 89516 19612
rect 89540 19610 89596 19612
rect 89300 19558 89346 19610
rect 89346 19558 89356 19610
rect 89380 19558 89410 19610
rect 89410 19558 89422 19610
rect 89422 19558 89436 19610
rect 89460 19558 89474 19610
rect 89474 19558 89486 19610
rect 89486 19558 89516 19610
rect 89540 19558 89550 19610
rect 89550 19558 89596 19610
rect 89300 19556 89356 19558
rect 89380 19556 89436 19558
rect 89460 19556 89516 19558
rect 89540 19556 89596 19558
rect 89300 18522 89356 18524
rect 89380 18522 89436 18524
rect 89460 18522 89516 18524
rect 89540 18522 89596 18524
rect 89300 18470 89346 18522
rect 89346 18470 89356 18522
rect 89380 18470 89410 18522
rect 89410 18470 89422 18522
rect 89422 18470 89436 18522
rect 89460 18470 89474 18522
rect 89474 18470 89486 18522
rect 89486 18470 89516 18522
rect 89540 18470 89550 18522
rect 89550 18470 89596 18522
rect 89300 18468 89356 18470
rect 89380 18468 89436 18470
rect 89460 18468 89516 18470
rect 89540 18468 89596 18470
rect 89300 17434 89356 17436
rect 89380 17434 89436 17436
rect 89460 17434 89516 17436
rect 89540 17434 89596 17436
rect 89300 17382 89346 17434
rect 89346 17382 89356 17434
rect 89380 17382 89410 17434
rect 89410 17382 89422 17434
rect 89422 17382 89436 17434
rect 89460 17382 89474 17434
rect 89474 17382 89486 17434
rect 89486 17382 89516 17434
rect 89540 17382 89550 17434
rect 89550 17382 89596 17434
rect 89300 17380 89356 17382
rect 89380 17380 89436 17382
rect 89460 17380 89516 17382
rect 89540 17380 89596 17382
rect 89300 16346 89356 16348
rect 89380 16346 89436 16348
rect 89460 16346 89516 16348
rect 89540 16346 89596 16348
rect 89300 16294 89346 16346
rect 89346 16294 89356 16346
rect 89380 16294 89410 16346
rect 89410 16294 89422 16346
rect 89422 16294 89436 16346
rect 89460 16294 89474 16346
rect 89474 16294 89486 16346
rect 89486 16294 89516 16346
rect 89540 16294 89550 16346
rect 89550 16294 89596 16346
rect 89300 16292 89356 16294
rect 89380 16292 89436 16294
rect 89460 16292 89516 16294
rect 89540 16292 89596 16294
rect 89300 15258 89356 15260
rect 89380 15258 89436 15260
rect 89460 15258 89516 15260
rect 89540 15258 89596 15260
rect 89300 15206 89346 15258
rect 89346 15206 89356 15258
rect 89380 15206 89410 15258
rect 89410 15206 89422 15258
rect 89422 15206 89436 15258
rect 89460 15206 89474 15258
rect 89474 15206 89486 15258
rect 89486 15206 89516 15258
rect 89540 15206 89550 15258
rect 89550 15206 89596 15258
rect 89300 15204 89356 15206
rect 89380 15204 89436 15206
rect 89460 15204 89516 15206
rect 89540 15204 89596 15206
rect 89300 14170 89356 14172
rect 89380 14170 89436 14172
rect 89460 14170 89516 14172
rect 89540 14170 89596 14172
rect 89300 14118 89346 14170
rect 89346 14118 89356 14170
rect 89380 14118 89410 14170
rect 89410 14118 89422 14170
rect 89422 14118 89436 14170
rect 89460 14118 89474 14170
rect 89474 14118 89486 14170
rect 89486 14118 89516 14170
rect 89540 14118 89550 14170
rect 89550 14118 89596 14170
rect 89300 14116 89356 14118
rect 89380 14116 89436 14118
rect 89460 14116 89516 14118
rect 89540 14116 89596 14118
rect 89300 13082 89356 13084
rect 89380 13082 89436 13084
rect 89460 13082 89516 13084
rect 89540 13082 89596 13084
rect 89300 13030 89346 13082
rect 89346 13030 89356 13082
rect 89380 13030 89410 13082
rect 89410 13030 89422 13082
rect 89422 13030 89436 13082
rect 89460 13030 89474 13082
rect 89474 13030 89486 13082
rect 89486 13030 89516 13082
rect 89540 13030 89550 13082
rect 89550 13030 89596 13082
rect 89300 13028 89356 13030
rect 89380 13028 89436 13030
rect 89460 13028 89516 13030
rect 89540 13028 89596 13030
rect 89300 11994 89356 11996
rect 89380 11994 89436 11996
rect 89460 11994 89516 11996
rect 89540 11994 89596 11996
rect 89300 11942 89346 11994
rect 89346 11942 89356 11994
rect 89380 11942 89410 11994
rect 89410 11942 89422 11994
rect 89422 11942 89436 11994
rect 89460 11942 89474 11994
rect 89474 11942 89486 11994
rect 89486 11942 89516 11994
rect 89540 11942 89550 11994
rect 89550 11942 89596 11994
rect 89300 11940 89356 11942
rect 89380 11940 89436 11942
rect 89460 11940 89516 11942
rect 89540 11940 89596 11942
rect 89300 10906 89356 10908
rect 89380 10906 89436 10908
rect 89460 10906 89516 10908
rect 89540 10906 89596 10908
rect 89300 10854 89346 10906
rect 89346 10854 89356 10906
rect 89380 10854 89410 10906
rect 89410 10854 89422 10906
rect 89422 10854 89436 10906
rect 89460 10854 89474 10906
rect 89474 10854 89486 10906
rect 89486 10854 89516 10906
rect 89540 10854 89550 10906
rect 89550 10854 89596 10906
rect 89300 10852 89356 10854
rect 89380 10852 89436 10854
rect 89460 10852 89516 10854
rect 89540 10852 89596 10854
rect 89300 9818 89356 9820
rect 89380 9818 89436 9820
rect 89460 9818 89516 9820
rect 89540 9818 89596 9820
rect 89300 9766 89346 9818
rect 89346 9766 89356 9818
rect 89380 9766 89410 9818
rect 89410 9766 89422 9818
rect 89422 9766 89436 9818
rect 89460 9766 89474 9818
rect 89474 9766 89486 9818
rect 89486 9766 89516 9818
rect 89540 9766 89550 9818
rect 89550 9766 89596 9818
rect 89300 9764 89356 9766
rect 89380 9764 89436 9766
rect 89460 9764 89516 9766
rect 89540 9764 89596 9766
rect 89300 8730 89356 8732
rect 89380 8730 89436 8732
rect 89460 8730 89516 8732
rect 89540 8730 89596 8732
rect 89300 8678 89346 8730
rect 89346 8678 89356 8730
rect 89380 8678 89410 8730
rect 89410 8678 89422 8730
rect 89422 8678 89436 8730
rect 89460 8678 89474 8730
rect 89474 8678 89486 8730
rect 89486 8678 89516 8730
rect 89540 8678 89550 8730
rect 89550 8678 89596 8730
rect 89300 8676 89356 8678
rect 89380 8676 89436 8678
rect 89460 8676 89516 8678
rect 89540 8676 89596 8678
rect 89300 7642 89356 7644
rect 89380 7642 89436 7644
rect 89460 7642 89516 7644
rect 89540 7642 89596 7644
rect 89300 7590 89346 7642
rect 89346 7590 89356 7642
rect 89380 7590 89410 7642
rect 89410 7590 89422 7642
rect 89422 7590 89436 7642
rect 89460 7590 89474 7642
rect 89474 7590 89486 7642
rect 89486 7590 89516 7642
rect 89540 7590 89550 7642
rect 89550 7590 89596 7642
rect 89300 7588 89356 7590
rect 89380 7588 89436 7590
rect 89460 7588 89516 7590
rect 89540 7588 89596 7590
rect 89300 6554 89356 6556
rect 89380 6554 89436 6556
rect 89460 6554 89516 6556
rect 89540 6554 89596 6556
rect 89300 6502 89346 6554
rect 89346 6502 89356 6554
rect 89380 6502 89410 6554
rect 89410 6502 89422 6554
rect 89422 6502 89436 6554
rect 89460 6502 89474 6554
rect 89474 6502 89486 6554
rect 89486 6502 89516 6554
rect 89540 6502 89550 6554
rect 89550 6502 89596 6554
rect 89300 6500 89356 6502
rect 89380 6500 89436 6502
rect 89460 6500 89516 6502
rect 89540 6500 89596 6502
rect 89300 5466 89356 5468
rect 89380 5466 89436 5468
rect 89460 5466 89516 5468
rect 89540 5466 89596 5468
rect 89300 5414 89346 5466
rect 89346 5414 89356 5466
rect 89380 5414 89410 5466
rect 89410 5414 89422 5466
rect 89422 5414 89436 5466
rect 89460 5414 89474 5466
rect 89474 5414 89486 5466
rect 89486 5414 89516 5466
rect 89540 5414 89550 5466
rect 89550 5414 89596 5466
rect 89300 5412 89356 5414
rect 89380 5412 89436 5414
rect 89460 5412 89516 5414
rect 89540 5412 89596 5414
rect 89300 4378 89356 4380
rect 89380 4378 89436 4380
rect 89460 4378 89516 4380
rect 89540 4378 89596 4380
rect 89300 4326 89346 4378
rect 89346 4326 89356 4378
rect 89380 4326 89410 4378
rect 89410 4326 89422 4378
rect 89422 4326 89436 4378
rect 89460 4326 89474 4378
rect 89474 4326 89486 4378
rect 89486 4326 89516 4378
rect 89540 4326 89550 4378
rect 89550 4326 89596 4378
rect 89300 4324 89356 4326
rect 89380 4324 89436 4326
rect 89460 4324 89516 4326
rect 89540 4324 89596 4326
rect 89300 3290 89356 3292
rect 89380 3290 89436 3292
rect 89460 3290 89516 3292
rect 89540 3290 89596 3292
rect 89300 3238 89346 3290
rect 89346 3238 89356 3290
rect 89380 3238 89410 3290
rect 89410 3238 89422 3290
rect 89422 3238 89436 3290
rect 89460 3238 89474 3290
rect 89474 3238 89486 3290
rect 89486 3238 89516 3290
rect 89540 3238 89550 3290
rect 89550 3238 89596 3290
rect 89300 3236 89356 3238
rect 89380 3236 89436 3238
rect 89460 3236 89516 3238
rect 89540 3236 89596 3238
rect 89534 2508 89590 2544
rect 89534 2488 89536 2508
rect 89536 2488 89588 2508
rect 89588 2488 89590 2508
rect 88982 1400 89038 1456
rect 89300 2202 89356 2204
rect 89380 2202 89436 2204
rect 89460 2202 89516 2204
rect 89540 2202 89596 2204
rect 89300 2150 89346 2202
rect 89346 2150 89356 2202
rect 89380 2150 89410 2202
rect 89410 2150 89422 2202
rect 89422 2150 89436 2202
rect 89460 2150 89474 2202
rect 89474 2150 89486 2202
rect 89486 2150 89516 2202
rect 89540 2150 89550 2202
rect 89550 2150 89596 2202
rect 89300 2148 89356 2150
rect 89380 2148 89436 2150
rect 89460 2148 89516 2150
rect 89540 2148 89596 2150
rect 89718 2080 89774 2136
rect 89442 1808 89498 1864
rect 89350 1436 89352 1456
rect 89352 1436 89404 1456
rect 89404 1436 89406 1456
rect 89350 1400 89406 1436
rect 89626 1672 89682 1728
rect 89810 1808 89866 1864
rect 91742 26868 91744 26888
rect 91744 26868 91796 26888
rect 91796 26868 91798 26888
rect 91742 26832 91798 26868
rect 92202 27240 92258 27296
rect 92754 26560 92810 26616
rect 92846 26424 92902 26480
rect 92202 2488 92258 2544
rect 90914 1400 90970 1456
rect 92294 2080 92350 2136
rect 95882 27512 95938 27568
rect 96710 27512 96766 27568
rect 96250 27376 96306 27432
rect 96434 27240 96490 27296
rect 96710 27276 96712 27296
rect 96712 27276 96764 27296
rect 96764 27276 96766 27296
rect 96710 27240 96766 27276
rect 97170 27104 97226 27160
rect 95790 26560 95846 26616
rect 95974 26288 96030 26344
rect 104024 27770 104080 27772
rect 104104 27770 104160 27772
rect 104184 27770 104240 27772
rect 104264 27770 104320 27772
rect 104024 27718 104070 27770
rect 104070 27718 104080 27770
rect 104104 27718 104134 27770
rect 104134 27718 104146 27770
rect 104146 27718 104160 27770
rect 104184 27718 104198 27770
rect 104198 27718 104210 27770
rect 104210 27718 104240 27770
rect 104264 27718 104274 27770
rect 104274 27718 104320 27770
rect 104024 27716 104080 27718
rect 104104 27716 104160 27718
rect 104184 27716 104240 27718
rect 104264 27716 104320 27718
rect 100206 26852 100262 26888
rect 100206 26832 100208 26852
rect 100208 26832 100260 26852
rect 100260 26832 100262 26852
rect 104990 27396 105046 27432
rect 104990 27376 104992 27396
rect 104992 27376 105044 27396
rect 105044 27376 105046 27396
rect 105634 27276 105636 27296
rect 105636 27276 105688 27296
rect 105688 27276 105690 27296
rect 105634 27240 105690 27276
rect 104898 26968 104954 27024
rect 104024 26682 104080 26684
rect 104104 26682 104160 26684
rect 104184 26682 104240 26684
rect 104264 26682 104320 26684
rect 104024 26630 104070 26682
rect 104070 26630 104080 26682
rect 104104 26630 104134 26682
rect 104134 26630 104146 26682
rect 104146 26630 104160 26682
rect 104184 26630 104198 26682
rect 104198 26630 104210 26682
rect 104210 26630 104240 26682
rect 104264 26630 104274 26682
rect 104274 26630 104320 26682
rect 104024 26628 104080 26630
rect 104104 26628 104160 26630
rect 104184 26628 104240 26630
rect 104264 26628 104320 26630
rect 104806 26832 104862 26888
rect 104024 25594 104080 25596
rect 104104 25594 104160 25596
rect 104184 25594 104240 25596
rect 104264 25594 104320 25596
rect 104024 25542 104070 25594
rect 104070 25542 104080 25594
rect 104104 25542 104134 25594
rect 104134 25542 104146 25594
rect 104146 25542 104160 25594
rect 104184 25542 104198 25594
rect 104198 25542 104210 25594
rect 104210 25542 104240 25594
rect 104264 25542 104274 25594
rect 104274 25542 104320 25594
rect 104024 25540 104080 25542
rect 104104 25540 104160 25542
rect 104184 25540 104240 25542
rect 104264 25540 104320 25542
rect 104024 24506 104080 24508
rect 104104 24506 104160 24508
rect 104184 24506 104240 24508
rect 104264 24506 104320 24508
rect 104024 24454 104070 24506
rect 104070 24454 104080 24506
rect 104104 24454 104134 24506
rect 104134 24454 104146 24506
rect 104146 24454 104160 24506
rect 104184 24454 104198 24506
rect 104198 24454 104210 24506
rect 104210 24454 104240 24506
rect 104264 24454 104274 24506
rect 104274 24454 104320 24506
rect 104024 24452 104080 24454
rect 104104 24452 104160 24454
rect 104184 24452 104240 24454
rect 104264 24452 104320 24454
rect 104024 23418 104080 23420
rect 104104 23418 104160 23420
rect 104184 23418 104240 23420
rect 104264 23418 104320 23420
rect 104024 23366 104070 23418
rect 104070 23366 104080 23418
rect 104104 23366 104134 23418
rect 104134 23366 104146 23418
rect 104146 23366 104160 23418
rect 104184 23366 104198 23418
rect 104198 23366 104210 23418
rect 104210 23366 104240 23418
rect 104264 23366 104274 23418
rect 104274 23366 104320 23418
rect 104024 23364 104080 23366
rect 104104 23364 104160 23366
rect 104184 23364 104240 23366
rect 104264 23364 104320 23366
rect 104024 22330 104080 22332
rect 104104 22330 104160 22332
rect 104184 22330 104240 22332
rect 104264 22330 104320 22332
rect 104024 22278 104070 22330
rect 104070 22278 104080 22330
rect 104104 22278 104134 22330
rect 104134 22278 104146 22330
rect 104146 22278 104160 22330
rect 104184 22278 104198 22330
rect 104198 22278 104210 22330
rect 104210 22278 104240 22330
rect 104264 22278 104274 22330
rect 104274 22278 104320 22330
rect 104024 22276 104080 22278
rect 104104 22276 104160 22278
rect 104184 22276 104240 22278
rect 104264 22276 104320 22278
rect 104024 21242 104080 21244
rect 104104 21242 104160 21244
rect 104184 21242 104240 21244
rect 104264 21242 104320 21244
rect 104024 21190 104070 21242
rect 104070 21190 104080 21242
rect 104104 21190 104134 21242
rect 104134 21190 104146 21242
rect 104146 21190 104160 21242
rect 104184 21190 104198 21242
rect 104198 21190 104210 21242
rect 104210 21190 104240 21242
rect 104264 21190 104274 21242
rect 104274 21190 104320 21242
rect 104024 21188 104080 21190
rect 104104 21188 104160 21190
rect 104184 21188 104240 21190
rect 104264 21188 104320 21190
rect 104024 20154 104080 20156
rect 104104 20154 104160 20156
rect 104184 20154 104240 20156
rect 104264 20154 104320 20156
rect 104024 20102 104070 20154
rect 104070 20102 104080 20154
rect 104104 20102 104134 20154
rect 104134 20102 104146 20154
rect 104146 20102 104160 20154
rect 104184 20102 104198 20154
rect 104198 20102 104210 20154
rect 104210 20102 104240 20154
rect 104264 20102 104274 20154
rect 104274 20102 104320 20154
rect 104024 20100 104080 20102
rect 104104 20100 104160 20102
rect 104184 20100 104240 20102
rect 104264 20100 104320 20102
rect 104024 19066 104080 19068
rect 104104 19066 104160 19068
rect 104184 19066 104240 19068
rect 104264 19066 104320 19068
rect 104024 19014 104070 19066
rect 104070 19014 104080 19066
rect 104104 19014 104134 19066
rect 104134 19014 104146 19066
rect 104146 19014 104160 19066
rect 104184 19014 104198 19066
rect 104198 19014 104210 19066
rect 104210 19014 104240 19066
rect 104264 19014 104274 19066
rect 104274 19014 104320 19066
rect 104024 19012 104080 19014
rect 104104 19012 104160 19014
rect 104184 19012 104240 19014
rect 104264 19012 104320 19014
rect 104024 17978 104080 17980
rect 104104 17978 104160 17980
rect 104184 17978 104240 17980
rect 104264 17978 104320 17980
rect 104024 17926 104070 17978
rect 104070 17926 104080 17978
rect 104104 17926 104134 17978
rect 104134 17926 104146 17978
rect 104146 17926 104160 17978
rect 104184 17926 104198 17978
rect 104198 17926 104210 17978
rect 104210 17926 104240 17978
rect 104264 17926 104274 17978
rect 104274 17926 104320 17978
rect 104024 17924 104080 17926
rect 104104 17924 104160 17926
rect 104184 17924 104240 17926
rect 104264 17924 104320 17926
rect 104024 16890 104080 16892
rect 104104 16890 104160 16892
rect 104184 16890 104240 16892
rect 104264 16890 104320 16892
rect 104024 16838 104070 16890
rect 104070 16838 104080 16890
rect 104104 16838 104134 16890
rect 104134 16838 104146 16890
rect 104146 16838 104160 16890
rect 104184 16838 104198 16890
rect 104198 16838 104210 16890
rect 104210 16838 104240 16890
rect 104264 16838 104274 16890
rect 104274 16838 104320 16890
rect 104024 16836 104080 16838
rect 104104 16836 104160 16838
rect 104184 16836 104240 16838
rect 104264 16836 104320 16838
rect 104024 15802 104080 15804
rect 104104 15802 104160 15804
rect 104184 15802 104240 15804
rect 104264 15802 104320 15804
rect 104024 15750 104070 15802
rect 104070 15750 104080 15802
rect 104104 15750 104134 15802
rect 104134 15750 104146 15802
rect 104146 15750 104160 15802
rect 104184 15750 104198 15802
rect 104198 15750 104210 15802
rect 104210 15750 104240 15802
rect 104264 15750 104274 15802
rect 104274 15750 104320 15802
rect 104024 15748 104080 15750
rect 104104 15748 104160 15750
rect 104184 15748 104240 15750
rect 104264 15748 104320 15750
rect 104024 14714 104080 14716
rect 104104 14714 104160 14716
rect 104184 14714 104240 14716
rect 104264 14714 104320 14716
rect 104024 14662 104070 14714
rect 104070 14662 104080 14714
rect 104104 14662 104134 14714
rect 104134 14662 104146 14714
rect 104146 14662 104160 14714
rect 104184 14662 104198 14714
rect 104198 14662 104210 14714
rect 104210 14662 104240 14714
rect 104264 14662 104274 14714
rect 104274 14662 104320 14714
rect 104024 14660 104080 14662
rect 104104 14660 104160 14662
rect 104184 14660 104240 14662
rect 104264 14660 104320 14662
rect 104024 13626 104080 13628
rect 104104 13626 104160 13628
rect 104184 13626 104240 13628
rect 104264 13626 104320 13628
rect 104024 13574 104070 13626
rect 104070 13574 104080 13626
rect 104104 13574 104134 13626
rect 104134 13574 104146 13626
rect 104146 13574 104160 13626
rect 104184 13574 104198 13626
rect 104198 13574 104210 13626
rect 104210 13574 104240 13626
rect 104264 13574 104274 13626
rect 104274 13574 104320 13626
rect 104024 13572 104080 13574
rect 104104 13572 104160 13574
rect 104184 13572 104240 13574
rect 104264 13572 104320 13574
rect 104024 12538 104080 12540
rect 104104 12538 104160 12540
rect 104184 12538 104240 12540
rect 104264 12538 104320 12540
rect 104024 12486 104070 12538
rect 104070 12486 104080 12538
rect 104104 12486 104134 12538
rect 104134 12486 104146 12538
rect 104146 12486 104160 12538
rect 104184 12486 104198 12538
rect 104198 12486 104210 12538
rect 104210 12486 104240 12538
rect 104264 12486 104274 12538
rect 104274 12486 104320 12538
rect 104024 12484 104080 12486
rect 104104 12484 104160 12486
rect 104184 12484 104240 12486
rect 104264 12484 104320 12486
rect 104024 11450 104080 11452
rect 104104 11450 104160 11452
rect 104184 11450 104240 11452
rect 104264 11450 104320 11452
rect 104024 11398 104070 11450
rect 104070 11398 104080 11450
rect 104104 11398 104134 11450
rect 104134 11398 104146 11450
rect 104146 11398 104160 11450
rect 104184 11398 104198 11450
rect 104198 11398 104210 11450
rect 104210 11398 104240 11450
rect 104264 11398 104274 11450
rect 104274 11398 104320 11450
rect 104024 11396 104080 11398
rect 104104 11396 104160 11398
rect 104184 11396 104240 11398
rect 104264 11396 104320 11398
rect 104024 10362 104080 10364
rect 104104 10362 104160 10364
rect 104184 10362 104240 10364
rect 104264 10362 104320 10364
rect 104024 10310 104070 10362
rect 104070 10310 104080 10362
rect 104104 10310 104134 10362
rect 104134 10310 104146 10362
rect 104146 10310 104160 10362
rect 104184 10310 104198 10362
rect 104198 10310 104210 10362
rect 104210 10310 104240 10362
rect 104264 10310 104274 10362
rect 104274 10310 104320 10362
rect 104024 10308 104080 10310
rect 104104 10308 104160 10310
rect 104184 10308 104240 10310
rect 104264 10308 104320 10310
rect 104024 9274 104080 9276
rect 104104 9274 104160 9276
rect 104184 9274 104240 9276
rect 104264 9274 104320 9276
rect 104024 9222 104070 9274
rect 104070 9222 104080 9274
rect 104104 9222 104134 9274
rect 104134 9222 104146 9274
rect 104146 9222 104160 9274
rect 104184 9222 104198 9274
rect 104198 9222 104210 9274
rect 104210 9222 104240 9274
rect 104264 9222 104274 9274
rect 104274 9222 104320 9274
rect 104024 9220 104080 9222
rect 104104 9220 104160 9222
rect 104184 9220 104240 9222
rect 104264 9220 104320 9222
rect 104024 8186 104080 8188
rect 104104 8186 104160 8188
rect 104184 8186 104240 8188
rect 104264 8186 104320 8188
rect 104024 8134 104070 8186
rect 104070 8134 104080 8186
rect 104104 8134 104134 8186
rect 104134 8134 104146 8186
rect 104146 8134 104160 8186
rect 104184 8134 104198 8186
rect 104198 8134 104210 8186
rect 104210 8134 104240 8186
rect 104264 8134 104274 8186
rect 104274 8134 104320 8186
rect 104024 8132 104080 8134
rect 104104 8132 104160 8134
rect 104184 8132 104240 8134
rect 104264 8132 104320 8134
rect 104024 7098 104080 7100
rect 104104 7098 104160 7100
rect 104184 7098 104240 7100
rect 104264 7098 104320 7100
rect 104024 7046 104070 7098
rect 104070 7046 104080 7098
rect 104104 7046 104134 7098
rect 104134 7046 104146 7098
rect 104146 7046 104160 7098
rect 104184 7046 104198 7098
rect 104198 7046 104210 7098
rect 104210 7046 104240 7098
rect 104264 7046 104274 7098
rect 104274 7046 104320 7098
rect 104024 7044 104080 7046
rect 104104 7044 104160 7046
rect 104184 7044 104240 7046
rect 104264 7044 104320 7046
rect 104024 6010 104080 6012
rect 104104 6010 104160 6012
rect 104184 6010 104240 6012
rect 104264 6010 104320 6012
rect 104024 5958 104070 6010
rect 104070 5958 104080 6010
rect 104104 5958 104134 6010
rect 104134 5958 104146 6010
rect 104146 5958 104160 6010
rect 104184 5958 104198 6010
rect 104198 5958 104210 6010
rect 104210 5958 104240 6010
rect 104264 5958 104274 6010
rect 104274 5958 104320 6010
rect 104024 5956 104080 5958
rect 104104 5956 104160 5958
rect 104184 5956 104240 5958
rect 104264 5956 104320 5958
rect 104024 4922 104080 4924
rect 104104 4922 104160 4924
rect 104184 4922 104240 4924
rect 104264 4922 104320 4924
rect 104024 4870 104070 4922
rect 104070 4870 104080 4922
rect 104104 4870 104134 4922
rect 104134 4870 104146 4922
rect 104146 4870 104160 4922
rect 104184 4870 104198 4922
rect 104198 4870 104210 4922
rect 104210 4870 104240 4922
rect 104264 4870 104274 4922
rect 104274 4870 104320 4922
rect 104024 4868 104080 4870
rect 104104 4868 104160 4870
rect 104184 4868 104240 4870
rect 104264 4868 104320 4870
rect 104024 3834 104080 3836
rect 104104 3834 104160 3836
rect 104184 3834 104240 3836
rect 104264 3834 104320 3836
rect 104024 3782 104070 3834
rect 104070 3782 104080 3834
rect 104104 3782 104134 3834
rect 104134 3782 104146 3834
rect 104146 3782 104160 3834
rect 104184 3782 104198 3834
rect 104198 3782 104210 3834
rect 104210 3782 104240 3834
rect 104264 3782 104274 3834
rect 104274 3782 104320 3834
rect 104024 3780 104080 3782
rect 104104 3780 104160 3782
rect 104184 3780 104240 3782
rect 104264 3780 104320 3782
rect 104024 2746 104080 2748
rect 104104 2746 104160 2748
rect 104184 2746 104240 2748
rect 104264 2746 104320 2748
rect 104024 2694 104070 2746
rect 104070 2694 104080 2746
rect 104104 2694 104134 2746
rect 104134 2694 104146 2746
rect 104146 2694 104160 2746
rect 104184 2694 104198 2746
rect 104198 2694 104210 2746
rect 104210 2694 104240 2746
rect 104264 2694 104274 2746
rect 104274 2694 104320 2746
rect 104024 2692 104080 2694
rect 104104 2692 104160 2694
rect 104184 2692 104240 2694
rect 104264 2692 104320 2694
rect 117134 29144 117190 29200
rect 117042 27920 117098 27976
rect 117318 27240 117374 27296
rect 115386 8880 115442 8936
rect 117226 23160 117282 23216
rect 117318 21120 117374 21176
rect 117226 16360 117282 16416
rect 117962 26560 118018 26616
rect 117962 25200 118018 25256
rect 117962 24556 117964 24576
rect 117964 24556 118016 24576
rect 118016 24556 118018 24576
rect 117962 24520 118018 24556
rect 117962 22500 118018 22536
rect 117962 22480 117964 22500
rect 117964 22480 118016 22500
rect 118016 22480 118018 22500
rect 117962 20440 118018 20496
rect 117962 19760 118018 19816
rect 117870 18400 117926 18456
rect 117318 11636 117320 11656
rect 117320 11636 117372 11656
rect 117372 11636 117374 11656
rect 117318 11600 117374 11636
rect 115570 2352 115626 2408
rect 116398 2080 116454 2136
rect 117870 17720 117926 17776
rect 117870 14356 117872 14376
rect 117872 14356 117924 14376
rect 117924 14356 117926 14376
rect 117870 14320 117926 14356
rect 117870 13640 117926 13696
rect 118146 15680 118202 15736
rect 117962 12960 118018 13016
rect 117962 10920 118018 10976
rect 117962 9560 118018 9616
rect 117962 8200 118018 8256
rect 117962 6840 118018 6896
rect 117870 6160 117926 6216
rect 117962 4800 118018 4856
rect 117778 4120 117834 4176
rect 116674 1400 116730 1456
rect 117870 2760 117926 2816
rect 117778 40 117834 96
<< metal3 >>
rect 119200 29338 120000 29368
rect 117270 29278 120000 29338
rect 117129 29202 117195 29205
rect 117270 29202 117330 29278
rect 119200 29248 120000 29278
rect 117129 29200 117330 29202
rect 117129 29144 117134 29200
rect 117190 29144 117330 29200
rect 117129 29142 117330 29144
rect 117129 29139 117195 29142
rect 0 28658 800 28688
rect 1209 28658 1275 28661
rect 0 28656 1275 28658
rect 0 28600 1214 28656
rect 1270 28600 1275 28656
rect 0 28598 1275 28600
rect 0 28568 800 28598
rect 1209 28595 1275 28598
rect 0 27978 800 28008
rect 2773 27978 2839 27981
rect 0 27976 2839 27978
rect 0 27920 2778 27976
rect 2834 27920 2839 27976
rect 0 27918 2839 27920
rect 0 27888 800 27918
rect 2773 27915 2839 27918
rect 40217 27978 40283 27981
rect 74901 27978 74967 27981
rect 85205 27978 85271 27981
rect 40217 27976 48330 27978
rect 40217 27920 40222 27976
rect 40278 27920 48330 27976
rect 40217 27918 48330 27920
rect 40217 27915 40283 27918
rect 29269 27842 29335 27845
rect 38285 27842 38351 27845
rect 29269 27840 38351 27842
rect 29269 27784 29274 27840
rect 29330 27784 38290 27840
rect 38346 27784 38351 27840
rect 29269 27782 38351 27784
rect 29269 27779 29335 27782
rect 38285 27779 38351 27782
rect 15670 27776 15986 27777
rect 15670 27712 15676 27776
rect 15740 27712 15756 27776
rect 15820 27712 15836 27776
rect 15900 27712 15916 27776
rect 15980 27712 15986 27776
rect 15670 27711 15986 27712
rect 45118 27776 45434 27777
rect 45118 27712 45124 27776
rect 45188 27712 45204 27776
rect 45268 27712 45284 27776
rect 45348 27712 45364 27776
rect 45428 27712 45434 27776
rect 45118 27711 45434 27712
rect 21173 27706 21239 27709
rect 34053 27706 34119 27709
rect 21173 27704 34119 27706
rect 21173 27648 21178 27704
rect 21234 27648 34058 27704
rect 34114 27648 34119 27704
rect 21173 27646 34119 27648
rect 48270 27706 48330 27918
rect 74901 27976 85271 27978
rect 74901 27920 74906 27976
rect 74962 27920 85210 27976
rect 85266 27920 85271 27976
rect 74901 27918 85271 27920
rect 74901 27915 74967 27918
rect 85205 27915 85271 27918
rect 117037 27978 117103 27981
rect 119200 27978 120000 28008
rect 117037 27976 120000 27978
rect 117037 27920 117042 27976
rect 117098 27920 120000 27976
rect 117037 27918 120000 27920
rect 117037 27915 117103 27918
rect 119200 27888 120000 27918
rect 49049 27842 49115 27845
rect 57053 27842 57119 27845
rect 49049 27840 57119 27842
rect 49049 27784 49054 27840
rect 49110 27784 57058 27840
rect 57114 27784 57119 27840
rect 49049 27782 57119 27784
rect 49049 27779 49115 27782
rect 57053 27779 57119 27782
rect 69933 27842 69999 27845
rect 73797 27842 73863 27845
rect 69933 27840 73863 27842
rect 69933 27784 69938 27840
rect 69994 27784 73802 27840
rect 73858 27784 73863 27840
rect 69933 27782 73863 27784
rect 69933 27779 69999 27782
rect 73797 27779 73863 27782
rect 74566 27776 74882 27777
rect 74566 27712 74572 27776
rect 74636 27712 74652 27776
rect 74716 27712 74732 27776
rect 74796 27712 74812 27776
rect 74876 27712 74882 27776
rect 74566 27711 74882 27712
rect 104014 27776 104330 27777
rect 104014 27712 104020 27776
rect 104084 27712 104100 27776
rect 104164 27712 104180 27776
rect 104244 27712 104260 27776
rect 104324 27712 104330 27776
rect 104014 27711 104330 27712
rect 60641 27706 60707 27709
rect 48270 27704 60707 27706
rect 48270 27648 60646 27704
rect 60702 27648 60707 27704
rect 48270 27646 60707 27648
rect 21173 27643 21239 27646
rect 34053 27643 34119 27646
rect 60641 27643 60707 27646
rect 60825 27706 60891 27709
rect 74257 27706 74323 27709
rect 60825 27704 74323 27706
rect 60825 27648 60830 27704
rect 60886 27648 74262 27704
rect 74318 27648 74323 27704
rect 60825 27646 74323 27648
rect 60825 27643 60891 27646
rect 74257 27643 74323 27646
rect 75177 27706 75243 27709
rect 79409 27706 79475 27709
rect 75177 27704 79475 27706
rect 75177 27648 75182 27704
rect 75238 27648 79414 27704
rect 79470 27648 79475 27704
rect 75177 27646 79475 27648
rect 75177 27643 75243 27646
rect 79409 27643 79475 27646
rect 23657 27570 23723 27573
rect 31109 27570 31175 27573
rect 23657 27568 31175 27570
rect 23657 27512 23662 27568
rect 23718 27512 31114 27568
rect 31170 27512 31175 27568
rect 23657 27510 31175 27512
rect 23657 27507 23723 27510
rect 31109 27507 31175 27510
rect 31385 27570 31451 27573
rect 33041 27570 33107 27573
rect 40677 27570 40743 27573
rect 31385 27568 32874 27570
rect 31385 27512 31390 27568
rect 31446 27512 32874 27568
rect 31385 27510 32874 27512
rect 31385 27507 31451 27510
rect 23565 27434 23631 27437
rect 30465 27434 30531 27437
rect 23565 27432 30531 27434
rect 23565 27376 23570 27432
rect 23626 27376 30470 27432
rect 30526 27376 30531 27432
rect 23565 27374 30531 27376
rect 23565 27371 23631 27374
rect 30465 27371 30531 27374
rect 30649 27434 30715 27437
rect 32121 27434 32187 27437
rect 30649 27432 32187 27434
rect 30649 27376 30654 27432
rect 30710 27376 32126 27432
rect 32182 27376 32187 27432
rect 30649 27374 32187 27376
rect 32814 27434 32874 27510
rect 33041 27568 40743 27570
rect 33041 27512 33046 27568
rect 33102 27512 40682 27568
rect 40738 27512 40743 27568
rect 33041 27510 40743 27512
rect 33041 27507 33107 27510
rect 40677 27507 40743 27510
rect 43805 27570 43871 27573
rect 50245 27570 50311 27573
rect 43805 27568 50311 27570
rect 43805 27512 43810 27568
rect 43866 27512 50250 27568
rect 50306 27512 50311 27568
rect 43805 27510 50311 27512
rect 43805 27507 43871 27510
rect 50245 27507 50311 27510
rect 50429 27570 50495 27573
rect 51809 27570 51875 27573
rect 50429 27568 51875 27570
rect 50429 27512 50434 27568
rect 50490 27512 51814 27568
rect 51870 27512 51875 27568
rect 50429 27510 51875 27512
rect 50429 27507 50495 27510
rect 51809 27507 51875 27510
rect 53281 27570 53347 27573
rect 60917 27570 60983 27573
rect 53281 27568 60983 27570
rect 53281 27512 53286 27568
rect 53342 27512 60922 27568
rect 60978 27512 60983 27568
rect 53281 27510 60983 27512
rect 53281 27507 53347 27510
rect 60917 27507 60983 27510
rect 61745 27570 61811 27573
rect 95877 27570 95943 27573
rect 96705 27570 96771 27573
rect 61745 27568 95943 27570
rect 61745 27512 61750 27568
rect 61806 27512 95882 27568
rect 95938 27512 95943 27568
rect 61745 27510 95943 27512
rect 61745 27507 61811 27510
rect 95877 27507 95943 27510
rect 96064 27568 96771 27570
rect 96064 27512 96710 27568
rect 96766 27512 96771 27568
rect 96064 27510 96771 27512
rect 35341 27434 35407 27437
rect 32814 27432 35407 27434
rect 32814 27376 35346 27432
rect 35402 27376 35407 27432
rect 32814 27374 35407 27376
rect 30649 27371 30715 27374
rect 32121 27371 32187 27374
rect 35341 27371 35407 27374
rect 37917 27434 37983 27437
rect 79041 27434 79107 27437
rect 37917 27432 79107 27434
rect 37917 27376 37922 27432
rect 37978 27376 79046 27432
rect 79102 27376 79107 27432
rect 37917 27374 79107 27376
rect 37917 27371 37983 27374
rect 79041 27371 79107 27374
rect 89069 27434 89135 27437
rect 96064 27434 96124 27510
rect 96705 27507 96771 27510
rect 89069 27432 96124 27434
rect 89069 27376 89074 27432
rect 89130 27376 96124 27432
rect 89069 27374 96124 27376
rect 96245 27434 96311 27437
rect 104985 27434 105051 27437
rect 96245 27432 105051 27434
rect 96245 27376 96250 27432
rect 96306 27376 104990 27432
rect 105046 27376 105051 27432
rect 96245 27374 105051 27376
rect 89069 27371 89135 27374
rect 96245 27371 96311 27374
rect 104985 27371 105051 27374
rect 14457 27298 14523 27301
rect 16205 27298 16271 27301
rect 14457 27296 16271 27298
rect 14457 27240 14462 27296
rect 14518 27240 16210 27296
rect 16266 27240 16271 27296
rect 14457 27238 16271 27240
rect 14457 27235 14523 27238
rect 16205 27235 16271 27238
rect 20621 27298 20687 27301
rect 30097 27298 30163 27301
rect 20621 27296 30163 27298
rect 20621 27240 20626 27296
rect 20682 27240 30102 27296
rect 30158 27240 30163 27296
rect 20621 27238 30163 27240
rect 20621 27235 20687 27238
rect 30097 27235 30163 27238
rect 33593 27298 33659 27301
rect 50429 27298 50495 27301
rect 33593 27296 50495 27298
rect 33593 27240 33598 27296
rect 33654 27240 50434 27296
rect 50490 27240 50495 27296
rect 33593 27238 50495 27240
rect 33593 27235 33659 27238
rect 50429 27235 50495 27238
rect 50613 27298 50679 27301
rect 53005 27298 53071 27301
rect 50613 27296 53071 27298
rect 50613 27240 50618 27296
rect 50674 27240 53010 27296
rect 53066 27240 53071 27296
rect 50613 27238 53071 27240
rect 50613 27235 50679 27238
rect 53005 27235 53071 27238
rect 53189 27298 53255 27301
rect 54017 27298 54083 27301
rect 55305 27298 55371 27301
rect 53189 27296 55371 27298
rect 53189 27240 53194 27296
rect 53250 27240 54022 27296
rect 54078 27240 55310 27296
rect 55366 27240 55371 27296
rect 53189 27238 55371 27240
rect 53189 27235 53255 27238
rect 54017 27235 54083 27238
rect 55305 27235 55371 27238
rect 56409 27298 56475 27301
rect 57697 27298 57763 27301
rect 56409 27296 57763 27298
rect 56409 27240 56414 27296
rect 56470 27240 57702 27296
rect 57758 27240 57763 27296
rect 56409 27238 57763 27240
rect 56409 27235 56475 27238
rect 57697 27235 57763 27238
rect 60917 27298 60983 27301
rect 68369 27298 68435 27301
rect 72417 27298 72483 27301
rect 60917 27296 62498 27298
rect 60917 27240 60922 27296
rect 60978 27240 62498 27296
rect 60917 27238 62498 27240
rect 60917 27235 60983 27238
rect 30394 27232 30710 27233
rect 30394 27168 30400 27232
rect 30464 27168 30480 27232
rect 30544 27168 30560 27232
rect 30624 27168 30640 27232
rect 30704 27168 30710 27232
rect 30394 27167 30710 27168
rect 59842 27232 60158 27233
rect 59842 27168 59848 27232
rect 59912 27168 59928 27232
rect 59992 27168 60008 27232
rect 60072 27168 60088 27232
rect 60152 27168 60158 27232
rect 59842 27167 60158 27168
rect 21909 27162 21975 27165
rect 25129 27162 25195 27165
rect 30189 27162 30255 27165
rect 21909 27160 22110 27162
rect 21909 27104 21914 27160
rect 21970 27104 22110 27160
rect 21909 27102 22110 27104
rect 21909 27099 21975 27102
rect 15193 27026 15259 27029
rect 21909 27026 21975 27029
rect 15193 27024 21975 27026
rect 15193 26968 15198 27024
rect 15254 26968 21914 27024
rect 21970 26968 21975 27024
rect 15193 26966 21975 26968
rect 22050 27026 22110 27102
rect 25129 27160 30255 27162
rect 25129 27104 25134 27160
rect 25190 27104 30194 27160
rect 30250 27104 30255 27160
rect 25129 27102 30255 27104
rect 25129 27099 25195 27102
rect 30189 27099 30255 27102
rect 40309 27162 40375 27165
rect 41873 27162 41939 27165
rect 40309 27160 41939 27162
rect 40309 27104 40314 27160
rect 40370 27104 41878 27160
rect 41934 27104 41939 27160
rect 40309 27102 41939 27104
rect 40309 27099 40375 27102
rect 41873 27099 41939 27102
rect 45921 27162 45987 27165
rect 50889 27162 50955 27165
rect 45921 27160 50955 27162
rect 45921 27104 45926 27160
rect 45982 27104 50894 27160
rect 50950 27104 50955 27160
rect 45921 27102 50955 27104
rect 45921 27099 45987 27102
rect 50889 27099 50955 27102
rect 53097 27162 53163 27165
rect 59537 27162 59603 27165
rect 53097 27160 59603 27162
rect 53097 27104 53102 27160
rect 53158 27104 59542 27160
rect 59598 27104 59603 27160
rect 53097 27102 59603 27104
rect 53097 27099 53163 27102
rect 59537 27099 59603 27102
rect 60733 27162 60799 27165
rect 62297 27162 62363 27165
rect 60733 27160 62363 27162
rect 60733 27104 60738 27160
rect 60794 27104 62302 27160
rect 62358 27104 62363 27160
rect 60733 27102 62363 27104
rect 62438 27162 62498 27238
rect 68369 27296 72483 27298
rect 68369 27240 68374 27296
rect 68430 27240 72422 27296
rect 72478 27240 72483 27296
rect 68369 27238 72483 27240
rect 68369 27235 68435 27238
rect 72417 27235 72483 27238
rect 78581 27298 78647 27301
rect 80237 27298 80303 27301
rect 78581 27296 80303 27298
rect 78581 27240 78586 27296
rect 78642 27240 80242 27296
rect 80298 27240 80303 27296
rect 78581 27238 80303 27240
rect 78581 27235 78647 27238
rect 80237 27235 80303 27238
rect 84469 27298 84535 27301
rect 85205 27298 85271 27301
rect 84469 27296 85271 27298
rect 84469 27240 84474 27296
rect 84530 27240 85210 27296
rect 85266 27240 85271 27296
rect 84469 27238 85271 27240
rect 84469 27235 84535 27238
rect 85205 27235 85271 27238
rect 92197 27298 92263 27301
rect 96429 27298 96495 27301
rect 92197 27296 96495 27298
rect 92197 27240 92202 27296
rect 92258 27240 96434 27296
rect 96490 27240 96495 27296
rect 92197 27238 96495 27240
rect 92197 27235 92263 27238
rect 96429 27235 96495 27238
rect 96705 27298 96771 27301
rect 105629 27298 105695 27301
rect 96705 27296 105695 27298
rect 96705 27240 96710 27296
rect 96766 27240 105634 27296
rect 105690 27240 105695 27296
rect 96705 27238 105695 27240
rect 96705 27235 96771 27238
rect 105629 27235 105695 27238
rect 117313 27298 117379 27301
rect 119200 27298 120000 27328
rect 117313 27296 120000 27298
rect 117313 27240 117318 27296
rect 117374 27240 120000 27296
rect 117313 27238 120000 27240
rect 117313 27235 117379 27238
rect 89290 27232 89606 27233
rect 89290 27168 89296 27232
rect 89360 27168 89376 27232
rect 89440 27168 89456 27232
rect 89520 27168 89536 27232
rect 89600 27168 89606 27232
rect 119200 27208 120000 27238
rect 89290 27167 89606 27168
rect 74809 27162 74875 27165
rect 62438 27160 74875 27162
rect 62438 27104 74814 27160
rect 74870 27104 74875 27160
rect 62438 27102 74875 27104
rect 60733 27099 60799 27102
rect 62297 27099 62363 27102
rect 74809 27099 74875 27102
rect 76557 27162 76623 27165
rect 79317 27162 79383 27165
rect 76557 27160 79383 27162
rect 76557 27104 76562 27160
rect 76618 27104 79322 27160
rect 79378 27104 79383 27160
rect 76557 27102 79383 27104
rect 76557 27099 76623 27102
rect 79317 27099 79383 27102
rect 80329 27162 80395 27165
rect 87321 27162 87387 27165
rect 80329 27160 87387 27162
rect 80329 27104 80334 27160
rect 80390 27104 87326 27160
rect 87382 27104 87387 27160
rect 80329 27102 87387 27104
rect 80329 27099 80395 27102
rect 87321 27099 87387 27102
rect 90357 27162 90423 27165
rect 97165 27162 97231 27165
rect 90357 27160 97231 27162
rect 90357 27104 90362 27160
rect 90418 27104 97170 27160
rect 97226 27104 97231 27160
rect 90357 27102 97231 27104
rect 90357 27099 90423 27102
rect 97165 27099 97231 27102
rect 22461 27026 22527 27029
rect 22050 27024 22527 27026
rect 22050 26968 22466 27024
rect 22522 26968 22527 27024
rect 22050 26966 22527 26968
rect 15193 26963 15259 26966
rect 21909 26963 21975 26966
rect 22461 26963 22527 26966
rect 26785 27026 26851 27029
rect 31569 27026 31635 27029
rect 26785 27024 31635 27026
rect 26785 26968 26790 27024
rect 26846 26968 31574 27024
rect 31630 26968 31635 27024
rect 26785 26966 31635 26968
rect 26785 26963 26851 26966
rect 31569 26963 31635 26966
rect 34605 27026 34671 27029
rect 35249 27026 35315 27029
rect 104893 27026 104959 27029
rect 34605 27024 104959 27026
rect 34605 26968 34610 27024
rect 34666 26968 35254 27024
rect 35310 26968 104898 27024
rect 104954 26968 104959 27024
rect 34605 26966 104959 26968
rect 34605 26963 34671 26966
rect 35249 26963 35315 26966
rect 104893 26963 104959 26966
rect 20713 26890 20779 26893
rect 75545 26890 75611 26893
rect 80053 26890 80119 26893
rect 20713 26888 75194 26890
rect 20713 26832 20718 26888
rect 20774 26832 75194 26888
rect 20713 26830 75194 26832
rect 20713 26827 20779 26830
rect 19701 26754 19767 26757
rect 22369 26754 22435 26757
rect 19701 26752 22435 26754
rect 19701 26696 19706 26752
rect 19762 26696 22374 26752
rect 22430 26696 22435 26752
rect 19701 26694 22435 26696
rect 19701 26691 19767 26694
rect 22369 26691 22435 26694
rect 24117 26754 24183 26757
rect 27153 26754 27219 26757
rect 24117 26752 27219 26754
rect 24117 26696 24122 26752
rect 24178 26696 27158 26752
rect 27214 26696 27219 26752
rect 24117 26694 27219 26696
rect 24117 26691 24183 26694
rect 27153 26691 27219 26694
rect 29269 26754 29335 26757
rect 40953 26754 41019 26757
rect 29269 26752 41019 26754
rect 29269 26696 29274 26752
rect 29330 26696 40958 26752
rect 41014 26696 41019 26752
rect 29269 26694 41019 26696
rect 29269 26691 29335 26694
rect 40953 26691 41019 26694
rect 50613 26754 50679 26757
rect 51165 26754 51231 26757
rect 50613 26752 51231 26754
rect 50613 26696 50618 26752
rect 50674 26696 51170 26752
rect 51226 26696 51231 26752
rect 50613 26694 51231 26696
rect 50613 26691 50679 26694
rect 51165 26691 51231 26694
rect 57237 26754 57303 26757
rect 60365 26754 60431 26757
rect 57237 26752 60431 26754
rect 57237 26696 57242 26752
rect 57298 26696 60370 26752
rect 60426 26696 60431 26752
rect 57237 26694 60431 26696
rect 57237 26691 57303 26694
rect 60365 26691 60431 26694
rect 60549 26754 60615 26757
rect 62297 26754 62363 26757
rect 60549 26752 62363 26754
rect 60549 26696 60554 26752
rect 60610 26696 62302 26752
rect 62358 26696 62363 26752
rect 60549 26694 62363 26696
rect 60549 26691 60615 26694
rect 62297 26691 62363 26694
rect 62481 26754 62547 26757
rect 69565 26754 69631 26757
rect 62481 26752 69631 26754
rect 62481 26696 62486 26752
rect 62542 26696 69570 26752
rect 69626 26696 69631 26752
rect 62481 26694 69631 26696
rect 62481 26691 62547 26694
rect 69565 26691 69631 26694
rect 69841 26754 69907 26757
rect 70342 26754 70348 26756
rect 69841 26752 70348 26754
rect 69841 26696 69846 26752
rect 69902 26696 70348 26752
rect 69841 26694 70348 26696
rect 69841 26691 69907 26694
rect 70342 26692 70348 26694
rect 70412 26692 70418 26756
rect 70485 26754 70551 26757
rect 73061 26754 73127 26757
rect 70485 26752 73127 26754
rect 70485 26696 70490 26752
rect 70546 26696 73066 26752
rect 73122 26696 73127 26752
rect 70485 26694 73127 26696
rect 75134 26754 75194 26830
rect 75545 26888 80119 26890
rect 75545 26832 75550 26888
rect 75606 26832 80058 26888
rect 80114 26832 80119 26888
rect 75545 26830 80119 26832
rect 75545 26827 75611 26830
rect 80053 26827 80119 26830
rect 80237 26890 80303 26893
rect 91737 26890 91803 26893
rect 80237 26888 91803 26890
rect 80237 26832 80242 26888
rect 80298 26832 91742 26888
rect 91798 26832 91803 26888
rect 80237 26830 91803 26832
rect 80237 26827 80303 26830
rect 91737 26827 91803 26830
rect 100201 26890 100267 26893
rect 104801 26890 104867 26893
rect 100201 26888 104867 26890
rect 100201 26832 100206 26888
rect 100262 26832 104806 26888
rect 104862 26832 104867 26888
rect 100201 26830 104867 26832
rect 100201 26827 100267 26830
rect 104801 26827 104867 26830
rect 81157 26754 81223 26757
rect 75134 26752 81223 26754
rect 75134 26696 81162 26752
rect 81218 26696 81223 26752
rect 75134 26694 81223 26696
rect 70485 26691 70551 26694
rect 73061 26691 73127 26694
rect 81157 26691 81223 26694
rect 15670 26688 15986 26689
rect 0 26618 800 26648
rect 15670 26624 15676 26688
rect 15740 26624 15756 26688
rect 15820 26624 15836 26688
rect 15900 26624 15916 26688
rect 15980 26624 15986 26688
rect 15670 26623 15986 26624
rect 45118 26688 45434 26689
rect 45118 26624 45124 26688
rect 45188 26624 45204 26688
rect 45268 26624 45284 26688
rect 45348 26624 45364 26688
rect 45428 26624 45434 26688
rect 45118 26623 45434 26624
rect 74566 26688 74882 26689
rect 74566 26624 74572 26688
rect 74636 26624 74652 26688
rect 74716 26624 74732 26688
rect 74796 26624 74812 26688
rect 74876 26624 74882 26688
rect 74566 26623 74882 26624
rect 104014 26688 104330 26689
rect 104014 26624 104020 26688
rect 104084 26624 104100 26688
rect 104164 26624 104180 26688
rect 104244 26624 104260 26688
rect 104324 26624 104330 26688
rect 104014 26623 104330 26624
rect 1393 26618 1459 26621
rect 0 26616 1459 26618
rect 0 26560 1398 26616
rect 1454 26560 1459 26616
rect 0 26558 1459 26560
rect 0 26528 800 26558
rect 1393 26555 1459 26558
rect 22461 26618 22527 26621
rect 31477 26618 31543 26621
rect 22461 26616 31543 26618
rect 22461 26560 22466 26616
rect 22522 26560 31482 26616
rect 31538 26560 31543 26616
rect 22461 26558 31543 26560
rect 22461 26555 22527 26558
rect 31477 26555 31543 26558
rect 33593 26618 33659 26621
rect 34973 26618 35039 26621
rect 33593 26616 35039 26618
rect 33593 26560 33598 26616
rect 33654 26560 34978 26616
rect 35034 26560 35039 26616
rect 33593 26558 35039 26560
rect 33593 26555 33659 26558
rect 34973 26555 35039 26558
rect 35157 26618 35223 26621
rect 38377 26618 38443 26621
rect 35157 26616 38443 26618
rect 35157 26560 35162 26616
rect 35218 26560 38382 26616
rect 38438 26560 38443 26616
rect 35157 26558 38443 26560
rect 35157 26555 35223 26558
rect 38377 26555 38443 26558
rect 41137 26618 41203 26621
rect 44081 26618 44147 26621
rect 41137 26616 44147 26618
rect 41137 26560 41142 26616
rect 41198 26560 44086 26616
rect 44142 26560 44147 26616
rect 41137 26558 44147 26560
rect 41137 26555 41203 26558
rect 44081 26555 44147 26558
rect 50521 26618 50587 26621
rect 51257 26618 51323 26621
rect 59169 26618 59235 26621
rect 50521 26616 51323 26618
rect 50521 26560 50526 26616
rect 50582 26560 51262 26616
rect 51318 26560 51323 26616
rect 50521 26558 51323 26560
rect 50521 26555 50587 26558
rect 51257 26555 51323 26558
rect 51398 26616 59235 26618
rect 51398 26560 59174 26616
rect 59230 26560 59235 26616
rect 51398 26558 59235 26560
rect 20345 26482 20411 26485
rect 28165 26482 28231 26485
rect 20345 26480 28231 26482
rect 20345 26424 20350 26480
rect 20406 26424 28170 26480
rect 28226 26424 28231 26480
rect 20345 26422 28231 26424
rect 20345 26419 20411 26422
rect 28165 26419 28231 26422
rect 28993 26482 29059 26485
rect 33869 26482 33935 26485
rect 28993 26480 33935 26482
rect 28993 26424 28998 26480
rect 29054 26424 33874 26480
rect 33930 26424 33935 26480
rect 28993 26422 33935 26424
rect 28993 26419 29059 26422
rect 33869 26419 33935 26422
rect 35801 26482 35867 26485
rect 38561 26482 38627 26485
rect 35801 26480 38627 26482
rect 35801 26424 35806 26480
rect 35862 26424 38566 26480
rect 38622 26424 38627 26480
rect 35801 26422 38627 26424
rect 35801 26419 35867 26422
rect 38561 26419 38627 26422
rect 40953 26482 41019 26485
rect 43437 26482 43503 26485
rect 50153 26482 50219 26485
rect 40953 26480 41430 26482
rect 40953 26424 40958 26480
rect 41014 26424 41430 26480
rect 40953 26422 41430 26424
rect 40953 26419 41019 26422
rect 22369 26346 22435 26349
rect 24485 26346 24551 26349
rect 22369 26344 24551 26346
rect 22369 26288 22374 26344
rect 22430 26288 24490 26344
rect 24546 26288 24551 26344
rect 22369 26286 24551 26288
rect 22369 26283 22435 26286
rect 24485 26283 24551 26286
rect 31569 26346 31635 26349
rect 31845 26346 31911 26349
rect 31569 26344 31911 26346
rect 31569 26288 31574 26344
rect 31630 26288 31850 26344
rect 31906 26288 31911 26344
rect 31569 26286 31911 26288
rect 31569 26283 31635 26286
rect 31845 26283 31911 26286
rect 32029 26346 32095 26349
rect 41229 26346 41295 26349
rect 32029 26344 41295 26346
rect 32029 26288 32034 26344
rect 32090 26288 41234 26344
rect 41290 26288 41295 26344
rect 32029 26286 41295 26288
rect 32029 26283 32095 26286
rect 41229 26283 41295 26286
rect 41370 26210 41430 26422
rect 43437 26480 50219 26482
rect 43437 26424 43442 26480
rect 43498 26424 50158 26480
rect 50214 26424 50219 26480
rect 43437 26422 50219 26424
rect 43437 26419 43503 26422
rect 50153 26419 50219 26422
rect 50705 26482 50771 26485
rect 51398 26482 51458 26558
rect 59169 26555 59235 26558
rect 59721 26618 59787 26621
rect 60917 26618 60983 26621
rect 72233 26618 72299 26621
rect 59721 26616 60750 26618
rect 59721 26560 59726 26616
rect 59782 26560 60750 26616
rect 59721 26558 60750 26560
rect 59721 26555 59787 26558
rect 50705 26480 51458 26482
rect 50705 26424 50710 26480
rect 50766 26424 51458 26480
rect 50705 26422 51458 26424
rect 51809 26482 51875 26485
rect 60549 26482 60615 26485
rect 51809 26480 60615 26482
rect 51809 26424 51814 26480
rect 51870 26424 60554 26480
rect 60610 26424 60615 26480
rect 51809 26422 60615 26424
rect 60690 26482 60750 26558
rect 60917 26616 72299 26618
rect 60917 26560 60922 26616
rect 60978 26560 72238 26616
rect 72294 26560 72299 26616
rect 60917 26558 72299 26560
rect 60917 26555 60983 26558
rect 72233 26555 72299 26558
rect 78765 26618 78831 26621
rect 81893 26618 81959 26621
rect 78765 26616 81959 26618
rect 78765 26560 78770 26616
rect 78826 26560 81898 26616
rect 81954 26560 81959 26616
rect 78765 26558 81959 26560
rect 78765 26555 78831 26558
rect 81893 26555 81959 26558
rect 92749 26618 92815 26621
rect 95785 26618 95851 26621
rect 92749 26616 95851 26618
rect 92749 26560 92754 26616
rect 92810 26560 95790 26616
rect 95846 26560 95851 26616
rect 92749 26558 95851 26560
rect 92749 26555 92815 26558
rect 95785 26555 95851 26558
rect 117957 26618 118023 26621
rect 119200 26618 120000 26648
rect 117957 26616 120000 26618
rect 117957 26560 117962 26616
rect 118018 26560 120000 26616
rect 117957 26558 120000 26560
rect 117957 26555 118023 26558
rect 119200 26528 120000 26558
rect 61193 26482 61259 26485
rect 60690 26480 61259 26482
rect 60690 26424 61198 26480
rect 61254 26424 61259 26480
rect 60690 26422 61259 26424
rect 50705 26419 50771 26422
rect 51809 26419 51875 26422
rect 60549 26419 60615 26422
rect 61193 26419 61259 26422
rect 61745 26482 61811 26485
rect 65057 26482 65123 26485
rect 79685 26482 79751 26485
rect 81433 26482 81499 26485
rect 61745 26480 81499 26482
rect 61745 26424 61750 26480
rect 61806 26424 65062 26480
rect 65118 26424 79690 26480
rect 79746 26424 81438 26480
rect 81494 26424 81499 26480
rect 61745 26422 81499 26424
rect 61745 26419 61811 26422
rect 65057 26419 65123 26422
rect 79685 26419 79751 26422
rect 81433 26419 81499 26422
rect 89069 26482 89135 26485
rect 92841 26482 92907 26485
rect 89069 26480 92907 26482
rect 89069 26424 89074 26480
rect 89130 26424 92846 26480
rect 92902 26424 92907 26480
rect 89069 26422 92907 26424
rect 89069 26419 89135 26422
rect 92841 26419 92907 26422
rect 41781 26346 41847 26349
rect 50153 26346 50219 26349
rect 41781 26344 50219 26346
rect 41781 26288 41786 26344
rect 41842 26288 50158 26344
rect 50214 26288 50219 26344
rect 41781 26286 50219 26288
rect 41781 26283 41847 26286
rect 50153 26283 50219 26286
rect 50981 26346 51047 26349
rect 58433 26346 58499 26349
rect 50981 26344 58499 26346
rect 50981 26288 50986 26344
rect 51042 26288 58438 26344
rect 58494 26288 58499 26344
rect 50981 26286 58499 26288
rect 50981 26283 51047 26286
rect 58433 26283 58499 26286
rect 60641 26346 60707 26349
rect 62205 26346 62271 26349
rect 60641 26344 62271 26346
rect 60641 26288 60646 26344
rect 60702 26288 62210 26344
rect 62266 26288 62271 26344
rect 60641 26286 62271 26288
rect 60641 26283 60707 26286
rect 62205 26283 62271 26286
rect 70710 26284 70716 26348
rect 70780 26346 70786 26348
rect 80237 26346 80303 26349
rect 70780 26344 80303 26346
rect 70780 26288 80242 26344
rect 80298 26288 80303 26344
rect 70780 26286 80303 26288
rect 70780 26284 70786 26286
rect 80237 26283 80303 26286
rect 80421 26346 80487 26349
rect 95969 26346 96035 26349
rect 80421 26344 96035 26346
rect 80421 26288 80426 26344
rect 80482 26288 95974 26344
rect 96030 26288 96035 26344
rect 80421 26286 96035 26288
rect 80421 26283 80487 26286
rect 95969 26283 96035 26286
rect 47117 26210 47183 26213
rect 41370 26208 47183 26210
rect 41370 26152 47122 26208
rect 47178 26152 47183 26208
rect 41370 26150 47183 26152
rect 47117 26147 47183 26150
rect 50889 26210 50955 26213
rect 51625 26210 51691 26213
rect 50889 26208 51691 26210
rect 50889 26152 50894 26208
rect 50950 26152 51630 26208
rect 51686 26152 51691 26208
rect 50889 26150 51691 26152
rect 50889 26147 50955 26150
rect 51625 26147 51691 26150
rect 63217 26210 63283 26213
rect 70485 26210 70551 26213
rect 63217 26208 70551 26210
rect 63217 26152 63222 26208
rect 63278 26152 70490 26208
rect 70546 26152 70551 26208
rect 63217 26150 70551 26152
rect 63217 26147 63283 26150
rect 70485 26147 70551 26150
rect 71865 26210 71931 26213
rect 79777 26210 79843 26213
rect 71865 26208 79843 26210
rect 71865 26152 71870 26208
rect 71926 26152 79782 26208
rect 79838 26152 79843 26208
rect 71865 26150 79843 26152
rect 71865 26147 71931 26150
rect 79777 26147 79843 26150
rect 30394 26144 30710 26145
rect 30394 26080 30400 26144
rect 30464 26080 30480 26144
rect 30544 26080 30560 26144
rect 30624 26080 30640 26144
rect 30704 26080 30710 26144
rect 30394 26079 30710 26080
rect 59842 26144 60158 26145
rect 59842 26080 59848 26144
rect 59912 26080 59928 26144
rect 59992 26080 60008 26144
rect 60072 26080 60088 26144
rect 60152 26080 60158 26144
rect 59842 26079 60158 26080
rect 89290 26144 89606 26145
rect 89290 26080 89296 26144
rect 89360 26080 89376 26144
rect 89440 26080 89456 26144
rect 89520 26080 89536 26144
rect 89600 26080 89606 26144
rect 89290 26079 89606 26080
rect 40769 26074 40835 26077
rect 47301 26074 47367 26077
rect 40769 26072 47367 26074
rect 40769 26016 40774 26072
rect 40830 26016 47306 26072
rect 47362 26016 47367 26072
rect 40769 26014 47367 26016
rect 40769 26011 40835 26014
rect 47301 26011 47367 26014
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 59629 25938 59695 25941
rect 69013 25938 69079 25941
rect 72509 25938 72575 25941
rect 59629 25936 72575 25938
rect 59629 25880 59634 25936
rect 59690 25880 69018 25936
rect 69074 25880 72514 25936
rect 72570 25880 72575 25936
rect 59629 25878 72575 25880
rect 59629 25875 59695 25878
rect 69013 25875 69079 25878
rect 72509 25875 72575 25878
rect 15670 25600 15986 25601
rect 15670 25536 15676 25600
rect 15740 25536 15756 25600
rect 15820 25536 15836 25600
rect 15900 25536 15916 25600
rect 15980 25536 15986 25600
rect 15670 25535 15986 25536
rect 45118 25600 45434 25601
rect 45118 25536 45124 25600
rect 45188 25536 45204 25600
rect 45268 25536 45284 25600
rect 45348 25536 45364 25600
rect 45428 25536 45434 25600
rect 45118 25535 45434 25536
rect 74566 25600 74882 25601
rect 74566 25536 74572 25600
rect 74636 25536 74652 25600
rect 74716 25536 74732 25600
rect 74796 25536 74812 25600
rect 74876 25536 74882 25600
rect 74566 25535 74882 25536
rect 104014 25600 104330 25601
rect 104014 25536 104020 25600
rect 104084 25536 104100 25600
rect 104164 25536 104180 25600
rect 104244 25536 104260 25600
rect 104324 25536 104330 25600
rect 104014 25535 104330 25536
rect 117957 25258 118023 25261
rect 119200 25258 120000 25288
rect 117957 25256 120000 25258
rect 117957 25200 117962 25256
rect 118018 25200 120000 25256
rect 117957 25198 120000 25200
rect 117957 25195 118023 25198
rect 119200 25168 120000 25198
rect 30394 25056 30710 25057
rect 30394 24992 30400 25056
rect 30464 24992 30480 25056
rect 30544 24992 30560 25056
rect 30624 24992 30640 25056
rect 30704 24992 30710 25056
rect 30394 24991 30710 24992
rect 59842 25056 60158 25057
rect 59842 24992 59848 25056
rect 59912 24992 59928 25056
rect 59992 24992 60008 25056
rect 60072 24992 60088 25056
rect 60152 24992 60158 25056
rect 59842 24991 60158 24992
rect 89290 25056 89606 25057
rect 89290 24992 89296 25056
rect 89360 24992 89376 25056
rect 89440 24992 89456 25056
rect 89520 24992 89536 25056
rect 89600 24992 89606 25056
rect 89290 24991 89606 24992
rect 0 24578 800 24608
rect 1393 24578 1459 24581
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 800 24518
rect 1393 24515 1459 24518
rect 117957 24578 118023 24581
rect 119200 24578 120000 24608
rect 117957 24576 120000 24578
rect 117957 24520 117962 24576
rect 118018 24520 120000 24576
rect 117957 24518 120000 24520
rect 117957 24515 118023 24518
rect 15670 24512 15986 24513
rect 15670 24448 15676 24512
rect 15740 24448 15756 24512
rect 15820 24448 15836 24512
rect 15900 24448 15916 24512
rect 15980 24448 15986 24512
rect 15670 24447 15986 24448
rect 45118 24512 45434 24513
rect 45118 24448 45124 24512
rect 45188 24448 45204 24512
rect 45268 24448 45284 24512
rect 45348 24448 45364 24512
rect 45428 24448 45434 24512
rect 45118 24447 45434 24448
rect 74566 24512 74882 24513
rect 74566 24448 74572 24512
rect 74636 24448 74652 24512
rect 74716 24448 74732 24512
rect 74796 24448 74812 24512
rect 74876 24448 74882 24512
rect 74566 24447 74882 24448
rect 104014 24512 104330 24513
rect 104014 24448 104020 24512
rect 104084 24448 104100 24512
rect 104164 24448 104180 24512
rect 104244 24448 104260 24512
rect 104324 24448 104330 24512
rect 119200 24488 120000 24518
rect 104014 24447 104330 24448
rect 30394 23968 30710 23969
rect 0 23898 800 23928
rect 30394 23904 30400 23968
rect 30464 23904 30480 23968
rect 30544 23904 30560 23968
rect 30624 23904 30640 23968
rect 30704 23904 30710 23968
rect 30394 23903 30710 23904
rect 59842 23968 60158 23969
rect 59842 23904 59848 23968
rect 59912 23904 59928 23968
rect 59992 23904 60008 23968
rect 60072 23904 60088 23968
rect 60152 23904 60158 23968
rect 59842 23903 60158 23904
rect 89290 23968 89606 23969
rect 89290 23904 89296 23968
rect 89360 23904 89376 23968
rect 89440 23904 89456 23968
rect 89520 23904 89536 23968
rect 89600 23904 89606 23968
rect 89290 23903 89606 23904
rect 1393 23898 1459 23901
rect 0 23896 1459 23898
rect 0 23840 1398 23896
rect 1454 23840 1459 23896
rect 0 23838 1459 23840
rect 0 23808 800 23838
rect 1393 23835 1459 23838
rect 15670 23424 15986 23425
rect 15670 23360 15676 23424
rect 15740 23360 15756 23424
rect 15820 23360 15836 23424
rect 15900 23360 15916 23424
rect 15980 23360 15986 23424
rect 15670 23359 15986 23360
rect 45118 23424 45434 23425
rect 45118 23360 45124 23424
rect 45188 23360 45204 23424
rect 45268 23360 45284 23424
rect 45348 23360 45364 23424
rect 45428 23360 45434 23424
rect 45118 23359 45434 23360
rect 74566 23424 74882 23425
rect 74566 23360 74572 23424
rect 74636 23360 74652 23424
rect 74716 23360 74732 23424
rect 74796 23360 74812 23424
rect 74876 23360 74882 23424
rect 74566 23359 74882 23360
rect 104014 23424 104330 23425
rect 104014 23360 104020 23424
rect 104084 23360 104100 23424
rect 104164 23360 104180 23424
rect 104244 23360 104260 23424
rect 104324 23360 104330 23424
rect 104014 23359 104330 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 117221 23218 117287 23221
rect 119200 23218 120000 23248
rect 117221 23216 120000 23218
rect 117221 23160 117226 23216
rect 117282 23160 120000 23216
rect 117221 23158 120000 23160
rect 117221 23155 117287 23158
rect 119200 23128 120000 23158
rect 30394 22880 30710 22881
rect 30394 22816 30400 22880
rect 30464 22816 30480 22880
rect 30544 22816 30560 22880
rect 30624 22816 30640 22880
rect 30704 22816 30710 22880
rect 30394 22815 30710 22816
rect 59842 22880 60158 22881
rect 59842 22816 59848 22880
rect 59912 22816 59928 22880
rect 59992 22816 60008 22880
rect 60072 22816 60088 22880
rect 60152 22816 60158 22880
rect 59842 22815 60158 22816
rect 89290 22880 89606 22881
rect 89290 22816 89296 22880
rect 89360 22816 89376 22880
rect 89440 22816 89456 22880
rect 89520 22816 89536 22880
rect 89600 22816 89606 22880
rect 89290 22815 89606 22816
rect 117957 22538 118023 22541
rect 119200 22538 120000 22568
rect 117957 22536 120000 22538
rect 117957 22480 117962 22536
rect 118018 22480 120000 22536
rect 117957 22478 120000 22480
rect 117957 22475 118023 22478
rect 119200 22448 120000 22478
rect 15670 22336 15986 22337
rect 15670 22272 15676 22336
rect 15740 22272 15756 22336
rect 15820 22272 15836 22336
rect 15900 22272 15916 22336
rect 15980 22272 15986 22336
rect 15670 22271 15986 22272
rect 45118 22336 45434 22337
rect 45118 22272 45124 22336
rect 45188 22272 45204 22336
rect 45268 22272 45284 22336
rect 45348 22272 45364 22336
rect 45428 22272 45434 22336
rect 45118 22271 45434 22272
rect 74566 22336 74882 22337
rect 74566 22272 74572 22336
rect 74636 22272 74652 22336
rect 74716 22272 74732 22336
rect 74796 22272 74812 22336
rect 74876 22272 74882 22336
rect 74566 22271 74882 22272
rect 104014 22336 104330 22337
rect 104014 22272 104020 22336
rect 104084 22272 104100 22336
rect 104164 22272 104180 22336
rect 104244 22272 104260 22336
rect 104324 22272 104330 22336
rect 104014 22271 104330 22272
rect 0 21858 800 21888
rect 1393 21858 1459 21861
rect 0 21856 1459 21858
rect 0 21800 1398 21856
rect 1454 21800 1459 21856
rect 0 21798 1459 21800
rect 0 21768 800 21798
rect 1393 21795 1459 21798
rect 30394 21792 30710 21793
rect 30394 21728 30400 21792
rect 30464 21728 30480 21792
rect 30544 21728 30560 21792
rect 30624 21728 30640 21792
rect 30704 21728 30710 21792
rect 30394 21727 30710 21728
rect 59842 21792 60158 21793
rect 59842 21728 59848 21792
rect 59912 21728 59928 21792
rect 59992 21728 60008 21792
rect 60072 21728 60088 21792
rect 60152 21728 60158 21792
rect 59842 21727 60158 21728
rect 89290 21792 89606 21793
rect 89290 21728 89296 21792
rect 89360 21728 89376 21792
rect 89440 21728 89456 21792
rect 89520 21728 89536 21792
rect 89600 21728 89606 21792
rect 89290 21727 89606 21728
rect 15670 21248 15986 21249
rect 0 21178 800 21208
rect 15670 21184 15676 21248
rect 15740 21184 15756 21248
rect 15820 21184 15836 21248
rect 15900 21184 15916 21248
rect 15980 21184 15986 21248
rect 15670 21183 15986 21184
rect 45118 21248 45434 21249
rect 45118 21184 45124 21248
rect 45188 21184 45204 21248
rect 45268 21184 45284 21248
rect 45348 21184 45364 21248
rect 45428 21184 45434 21248
rect 45118 21183 45434 21184
rect 74566 21248 74882 21249
rect 74566 21184 74572 21248
rect 74636 21184 74652 21248
rect 74716 21184 74732 21248
rect 74796 21184 74812 21248
rect 74876 21184 74882 21248
rect 74566 21183 74882 21184
rect 104014 21248 104330 21249
rect 104014 21184 104020 21248
rect 104084 21184 104100 21248
rect 104164 21184 104180 21248
rect 104244 21184 104260 21248
rect 104324 21184 104330 21248
rect 104014 21183 104330 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 800 21118
rect 1393 21115 1459 21118
rect 117313 21178 117379 21181
rect 119200 21178 120000 21208
rect 117313 21176 120000 21178
rect 117313 21120 117318 21176
rect 117374 21120 120000 21176
rect 117313 21118 120000 21120
rect 117313 21115 117379 21118
rect 119200 21088 120000 21118
rect 30394 20704 30710 20705
rect 30394 20640 30400 20704
rect 30464 20640 30480 20704
rect 30544 20640 30560 20704
rect 30624 20640 30640 20704
rect 30704 20640 30710 20704
rect 30394 20639 30710 20640
rect 59842 20704 60158 20705
rect 59842 20640 59848 20704
rect 59912 20640 59928 20704
rect 59992 20640 60008 20704
rect 60072 20640 60088 20704
rect 60152 20640 60158 20704
rect 59842 20639 60158 20640
rect 89290 20704 89606 20705
rect 89290 20640 89296 20704
rect 89360 20640 89376 20704
rect 89440 20640 89456 20704
rect 89520 20640 89536 20704
rect 89600 20640 89606 20704
rect 89290 20639 89606 20640
rect 117957 20498 118023 20501
rect 119200 20498 120000 20528
rect 117957 20496 120000 20498
rect 117957 20440 117962 20496
rect 118018 20440 120000 20496
rect 117957 20438 120000 20440
rect 117957 20435 118023 20438
rect 119200 20408 120000 20438
rect 15670 20160 15986 20161
rect 15670 20096 15676 20160
rect 15740 20096 15756 20160
rect 15820 20096 15836 20160
rect 15900 20096 15916 20160
rect 15980 20096 15986 20160
rect 15670 20095 15986 20096
rect 45118 20160 45434 20161
rect 45118 20096 45124 20160
rect 45188 20096 45204 20160
rect 45268 20096 45284 20160
rect 45348 20096 45364 20160
rect 45428 20096 45434 20160
rect 45118 20095 45434 20096
rect 74566 20160 74882 20161
rect 74566 20096 74572 20160
rect 74636 20096 74652 20160
rect 74716 20096 74732 20160
rect 74796 20096 74812 20160
rect 74876 20096 74882 20160
rect 74566 20095 74882 20096
rect 104014 20160 104330 20161
rect 104014 20096 104020 20160
rect 104084 20096 104100 20160
rect 104164 20096 104180 20160
rect 104244 20096 104260 20160
rect 104324 20096 104330 20160
rect 104014 20095 104330 20096
rect 0 19818 800 19848
rect 1393 19818 1459 19821
rect 0 19816 1459 19818
rect 0 19760 1398 19816
rect 1454 19760 1459 19816
rect 0 19758 1459 19760
rect 0 19728 800 19758
rect 1393 19755 1459 19758
rect 117957 19818 118023 19821
rect 119200 19818 120000 19848
rect 117957 19816 120000 19818
rect 117957 19760 117962 19816
rect 118018 19760 120000 19816
rect 117957 19758 120000 19760
rect 117957 19755 118023 19758
rect 119200 19728 120000 19758
rect 30394 19616 30710 19617
rect 30394 19552 30400 19616
rect 30464 19552 30480 19616
rect 30544 19552 30560 19616
rect 30624 19552 30640 19616
rect 30704 19552 30710 19616
rect 30394 19551 30710 19552
rect 59842 19616 60158 19617
rect 59842 19552 59848 19616
rect 59912 19552 59928 19616
rect 59992 19552 60008 19616
rect 60072 19552 60088 19616
rect 60152 19552 60158 19616
rect 59842 19551 60158 19552
rect 89290 19616 89606 19617
rect 89290 19552 89296 19616
rect 89360 19552 89376 19616
rect 89440 19552 89456 19616
rect 89520 19552 89536 19616
rect 89600 19552 89606 19616
rect 89290 19551 89606 19552
rect 0 19138 800 19168
rect 1853 19138 1919 19141
rect 0 19136 1919 19138
rect 0 19080 1858 19136
rect 1914 19080 1919 19136
rect 0 19078 1919 19080
rect 0 19048 800 19078
rect 1853 19075 1919 19078
rect 15670 19072 15986 19073
rect 15670 19008 15676 19072
rect 15740 19008 15756 19072
rect 15820 19008 15836 19072
rect 15900 19008 15916 19072
rect 15980 19008 15986 19072
rect 15670 19007 15986 19008
rect 45118 19072 45434 19073
rect 45118 19008 45124 19072
rect 45188 19008 45204 19072
rect 45268 19008 45284 19072
rect 45348 19008 45364 19072
rect 45428 19008 45434 19072
rect 45118 19007 45434 19008
rect 74566 19072 74882 19073
rect 74566 19008 74572 19072
rect 74636 19008 74652 19072
rect 74716 19008 74732 19072
rect 74796 19008 74812 19072
rect 74876 19008 74882 19072
rect 74566 19007 74882 19008
rect 104014 19072 104330 19073
rect 104014 19008 104020 19072
rect 104084 19008 104100 19072
rect 104164 19008 104180 19072
rect 104244 19008 104260 19072
rect 104324 19008 104330 19072
rect 104014 19007 104330 19008
rect 30394 18528 30710 18529
rect 0 18458 800 18488
rect 30394 18464 30400 18528
rect 30464 18464 30480 18528
rect 30544 18464 30560 18528
rect 30624 18464 30640 18528
rect 30704 18464 30710 18528
rect 30394 18463 30710 18464
rect 59842 18528 60158 18529
rect 59842 18464 59848 18528
rect 59912 18464 59928 18528
rect 59992 18464 60008 18528
rect 60072 18464 60088 18528
rect 60152 18464 60158 18528
rect 59842 18463 60158 18464
rect 89290 18528 89606 18529
rect 89290 18464 89296 18528
rect 89360 18464 89376 18528
rect 89440 18464 89456 18528
rect 89520 18464 89536 18528
rect 89600 18464 89606 18528
rect 89290 18463 89606 18464
rect 1393 18458 1459 18461
rect 0 18456 1459 18458
rect 0 18400 1398 18456
rect 1454 18400 1459 18456
rect 0 18398 1459 18400
rect 0 18368 800 18398
rect 1393 18395 1459 18398
rect 117865 18458 117931 18461
rect 119200 18458 120000 18488
rect 117865 18456 120000 18458
rect 117865 18400 117870 18456
rect 117926 18400 120000 18456
rect 117865 18398 120000 18400
rect 117865 18395 117931 18398
rect 119200 18368 120000 18398
rect 15670 17984 15986 17985
rect 15670 17920 15676 17984
rect 15740 17920 15756 17984
rect 15820 17920 15836 17984
rect 15900 17920 15916 17984
rect 15980 17920 15986 17984
rect 15670 17919 15986 17920
rect 45118 17984 45434 17985
rect 45118 17920 45124 17984
rect 45188 17920 45204 17984
rect 45268 17920 45284 17984
rect 45348 17920 45364 17984
rect 45428 17920 45434 17984
rect 45118 17919 45434 17920
rect 74566 17984 74882 17985
rect 74566 17920 74572 17984
rect 74636 17920 74652 17984
rect 74716 17920 74732 17984
rect 74796 17920 74812 17984
rect 74876 17920 74882 17984
rect 74566 17919 74882 17920
rect 104014 17984 104330 17985
rect 104014 17920 104020 17984
rect 104084 17920 104100 17984
rect 104164 17920 104180 17984
rect 104244 17920 104260 17984
rect 104324 17920 104330 17984
rect 104014 17919 104330 17920
rect 117865 17778 117931 17781
rect 119200 17778 120000 17808
rect 117865 17776 120000 17778
rect 117865 17720 117870 17776
rect 117926 17720 120000 17776
rect 117865 17718 120000 17720
rect 117865 17715 117931 17718
rect 119200 17688 120000 17718
rect 30394 17440 30710 17441
rect 30394 17376 30400 17440
rect 30464 17376 30480 17440
rect 30544 17376 30560 17440
rect 30624 17376 30640 17440
rect 30704 17376 30710 17440
rect 30394 17375 30710 17376
rect 59842 17440 60158 17441
rect 59842 17376 59848 17440
rect 59912 17376 59928 17440
rect 59992 17376 60008 17440
rect 60072 17376 60088 17440
rect 60152 17376 60158 17440
rect 59842 17375 60158 17376
rect 89290 17440 89606 17441
rect 89290 17376 89296 17440
rect 89360 17376 89376 17440
rect 89440 17376 89456 17440
rect 89520 17376 89536 17440
rect 89600 17376 89606 17440
rect 89290 17375 89606 17376
rect 0 17098 800 17128
rect 1393 17098 1459 17101
rect 0 17096 1459 17098
rect 0 17040 1398 17096
rect 1454 17040 1459 17096
rect 0 17038 1459 17040
rect 0 17008 800 17038
rect 1393 17035 1459 17038
rect 15670 16896 15986 16897
rect 15670 16832 15676 16896
rect 15740 16832 15756 16896
rect 15820 16832 15836 16896
rect 15900 16832 15916 16896
rect 15980 16832 15986 16896
rect 15670 16831 15986 16832
rect 45118 16896 45434 16897
rect 45118 16832 45124 16896
rect 45188 16832 45204 16896
rect 45268 16832 45284 16896
rect 45348 16832 45364 16896
rect 45428 16832 45434 16896
rect 45118 16831 45434 16832
rect 74566 16896 74882 16897
rect 74566 16832 74572 16896
rect 74636 16832 74652 16896
rect 74716 16832 74732 16896
rect 74796 16832 74812 16896
rect 74876 16832 74882 16896
rect 74566 16831 74882 16832
rect 104014 16896 104330 16897
rect 104014 16832 104020 16896
rect 104084 16832 104100 16896
rect 104164 16832 104180 16896
rect 104244 16832 104260 16896
rect 104324 16832 104330 16896
rect 104014 16831 104330 16832
rect 0 16418 800 16448
rect 1577 16418 1643 16421
rect 0 16416 1643 16418
rect 0 16360 1582 16416
rect 1638 16360 1643 16416
rect 0 16358 1643 16360
rect 0 16328 800 16358
rect 1577 16355 1643 16358
rect 117221 16418 117287 16421
rect 119200 16418 120000 16448
rect 117221 16416 120000 16418
rect 117221 16360 117226 16416
rect 117282 16360 120000 16416
rect 117221 16358 120000 16360
rect 117221 16355 117287 16358
rect 30394 16352 30710 16353
rect 30394 16288 30400 16352
rect 30464 16288 30480 16352
rect 30544 16288 30560 16352
rect 30624 16288 30640 16352
rect 30704 16288 30710 16352
rect 30394 16287 30710 16288
rect 59842 16352 60158 16353
rect 59842 16288 59848 16352
rect 59912 16288 59928 16352
rect 59992 16288 60008 16352
rect 60072 16288 60088 16352
rect 60152 16288 60158 16352
rect 59842 16287 60158 16288
rect 89290 16352 89606 16353
rect 89290 16288 89296 16352
rect 89360 16288 89376 16352
rect 89440 16288 89456 16352
rect 89520 16288 89536 16352
rect 89600 16288 89606 16352
rect 119200 16328 120000 16358
rect 89290 16287 89606 16288
rect 15670 15808 15986 15809
rect 15670 15744 15676 15808
rect 15740 15744 15756 15808
rect 15820 15744 15836 15808
rect 15900 15744 15916 15808
rect 15980 15744 15986 15808
rect 15670 15743 15986 15744
rect 45118 15808 45434 15809
rect 45118 15744 45124 15808
rect 45188 15744 45204 15808
rect 45268 15744 45284 15808
rect 45348 15744 45364 15808
rect 45428 15744 45434 15808
rect 45118 15743 45434 15744
rect 74566 15808 74882 15809
rect 74566 15744 74572 15808
rect 74636 15744 74652 15808
rect 74716 15744 74732 15808
rect 74796 15744 74812 15808
rect 74876 15744 74882 15808
rect 74566 15743 74882 15744
rect 104014 15808 104330 15809
rect 104014 15744 104020 15808
rect 104084 15744 104100 15808
rect 104164 15744 104180 15808
rect 104244 15744 104260 15808
rect 104324 15744 104330 15808
rect 104014 15743 104330 15744
rect 118141 15738 118207 15741
rect 119200 15738 120000 15768
rect 118141 15736 120000 15738
rect 118141 15680 118146 15736
rect 118202 15680 120000 15736
rect 118141 15678 120000 15680
rect 118141 15675 118207 15678
rect 119200 15648 120000 15678
rect 30394 15264 30710 15265
rect 30394 15200 30400 15264
rect 30464 15200 30480 15264
rect 30544 15200 30560 15264
rect 30624 15200 30640 15264
rect 30704 15200 30710 15264
rect 30394 15199 30710 15200
rect 59842 15264 60158 15265
rect 59842 15200 59848 15264
rect 59912 15200 59928 15264
rect 59992 15200 60008 15264
rect 60072 15200 60088 15264
rect 60152 15200 60158 15264
rect 59842 15199 60158 15200
rect 89290 15264 89606 15265
rect 89290 15200 89296 15264
rect 89360 15200 89376 15264
rect 89440 15200 89456 15264
rect 89520 15200 89536 15264
rect 89600 15200 89606 15264
rect 89290 15199 89606 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 68645 14922 68711 14925
rect 70209 14922 70275 14925
rect 68645 14920 70275 14922
rect 68645 14864 68650 14920
rect 68706 14864 70214 14920
rect 70270 14864 70275 14920
rect 68645 14862 70275 14864
rect 68645 14859 68711 14862
rect 70209 14859 70275 14862
rect 15670 14720 15986 14721
rect 15670 14656 15676 14720
rect 15740 14656 15756 14720
rect 15820 14656 15836 14720
rect 15900 14656 15916 14720
rect 15980 14656 15986 14720
rect 15670 14655 15986 14656
rect 45118 14720 45434 14721
rect 45118 14656 45124 14720
rect 45188 14656 45204 14720
rect 45268 14656 45284 14720
rect 45348 14656 45364 14720
rect 45428 14656 45434 14720
rect 45118 14655 45434 14656
rect 74566 14720 74882 14721
rect 74566 14656 74572 14720
rect 74636 14656 74652 14720
rect 74716 14656 74732 14720
rect 74796 14656 74812 14720
rect 74876 14656 74882 14720
rect 74566 14655 74882 14656
rect 104014 14720 104330 14721
rect 104014 14656 104020 14720
rect 104084 14656 104100 14720
rect 104164 14656 104180 14720
rect 104244 14656 104260 14720
rect 104324 14656 104330 14720
rect 104014 14655 104330 14656
rect 0 14378 800 14408
rect 1393 14378 1459 14381
rect 0 14376 1459 14378
rect 0 14320 1398 14376
rect 1454 14320 1459 14376
rect 0 14318 1459 14320
rect 0 14288 800 14318
rect 1393 14315 1459 14318
rect 117865 14378 117931 14381
rect 119200 14378 120000 14408
rect 117865 14376 120000 14378
rect 117865 14320 117870 14376
rect 117926 14320 120000 14376
rect 117865 14318 120000 14320
rect 117865 14315 117931 14318
rect 119200 14288 120000 14318
rect 30394 14176 30710 14177
rect 30394 14112 30400 14176
rect 30464 14112 30480 14176
rect 30544 14112 30560 14176
rect 30624 14112 30640 14176
rect 30704 14112 30710 14176
rect 30394 14111 30710 14112
rect 59842 14176 60158 14177
rect 59842 14112 59848 14176
rect 59912 14112 59928 14176
rect 59992 14112 60008 14176
rect 60072 14112 60088 14176
rect 60152 14112 60158 14176
rect 59842 14111 60158 14112
rect 89290 14176 89606 14177
rect 89290 14112 89296 14176
rect 89360 14112 89376 14176
rect 89440 14112 89456 14176
rect 89520 14112 89536 14176
rect 89600 14112 89606 14176
rect 89290 14111 89606 14112
rect 117865 13698 117931 13701
rect 119200 13698 120000 13728
rect 117865 13696 120000 13698
rect 117865 13640 117870 13696
rect 117926 13640 120000 13696
rect 117865 13638 120000 13640
rect 117865 13635 117931 13638
rect 15670 13632 15986 13633
rect 15670 13568 15676 13632
rect 15740 13568 15756 13632
rect 15820 13568 15836 13632
rect 15900 13568 15916 13632
rect 15980 13568 15986 13632
rect 15670 13567 15986 13568
rect 45118 13632 45434 13633
rect 45118 13568 45124 13632
rect 45188 13568 45204 13632
rect 45268 13568 45284 13632
rect 45348 13568 45364 13632
rect 45428 13568 45434 13632
rect 45118 13567 45434 13568
rect 74566 13632 74882 13633
rect 74566 13568 74572 13632
rect 74636 13568 74652 13632
rect 74716 13568 74732 13632
rect 74796 13568 74812 13632
rect 74876 13568 74882 13632
rect 74566 13567 74882 13568
rect 104014 13632 104330 13633
rect 104014 13568 104020 13632
rect 104084 13568 104100 13632
rect 104164 13568 104180 13632
rect 104244 13568 104260 13632
rect 104324 13568 104330 13632
rect 119200 13608 120000 13638
rect 104014 13567 104330 13568
rect 30394 13088 30710 13089
rect 0 13018 800 13048
rect 30394 13024 30400 13088
rect 30464 13024 30480 13088
rect 30544 13024 30560 13088
rect 30624 13024 30640 13088
rect 30704 13024 30710 13088
rect 30394 13023 30710 13024
rect 59842 13088 60158 13089
rect 59842 13024 59848 13088
rect 59912 13024 59928 13088
rect 59992 13024 60008 13088
rect 60072 13024 60088 13088
rect 60152 13024 60158 13088
rect 59842 13023 60158 13024
rect 89290 13088 89606 13089
rect 89290 13024 89296 13088
rect 89360 13024 89376 13088
rect 89440 13024 89456 13088
rect 89520 13024 89536 13088
rect 89600 13024 89606 13088
rect 89290 13023 89606 13024
rect 1853 13018 1919 13021
rect 0 13016 1919 13018
rect 0 12960 1858 13016
rect 1914 12960 1919 13016
rect 0 12958 1919 12960
rect 0 12928 800 12958
rect 1853 12955 1919 12958
rect 117957 13018 118023 13021
rect 119200 13018 120000 13048
rect 117957 13016 120000 13018
rect 117957 12960 117962 13016
rect 118018 12960 120000 13016
rect 117957 12958 120000 12960
rect 117957 12955 118023 12958
rect 119200 12928 120000 12958
rect 15670 12544 15986 12545
rect 15670 12480 15676 12544
rect 15740 12480 15756 12544
rect 15820 12480 15836 12544
rect 15900 12480 15916 12544
rect 15980 12480 15986 12544
rect 15670 12479 15986 12480
rect 45118 12544 45434 12545
rect 45118 12480 45124 12544
rect 45188 12480 45204 12544
rect 45268 12480 45284 12544
rect 45348 12480 45364 12544
rect 45428 12480 45434 12544
rect 45118 12479 45434 12480
rect 74566 12544 74882 12545
rect 74566 12480 74572 12544
rect 74636 12480 74652 12544
rect 74716 12480 74732 12544
rect 74796 12480 74812 12544
rect 74876 12480 74882 12544
rect 74566 12479 74882 12480
rect 104014 12544 104330 12545
rect 104014 12480 104020 12544
rect 104084 12480 104100 12544
rect 104164 12480 104180 12544
rect 104244 12480 104260 12544
rect 104324 12480 104330 12544
rect 104014 12479 104330 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 30394 12000 30710 12001
rect 30394 11936 30400 12000
rect 30464 11936 30480 12000
rect 30544 11936 30560 12000
rect 30624 11936 30640 12000
rect 30704 11936 30710 12000
rect 30394 11935 30710 11936
rect 59842 12000 60158 12001
rect 59842 11936 59848 12000
rect 59912 11936 59928 12000
rect 59992 11936 60008 12000
rect 60072 11936 60088 12000
rect 60152 11936 60158 12000
rect 59842 11935 60158 11936
rect 89290 12000 89606 12001
rect 89290 11936 89296 12000
rect 89360 11936 89376 12000
rect 89440 11936 89456 12000
rect 89520 11936 89536 12000
rect 89600 11936 89606 12000
rect 89290 11935 89606 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 117313 11658 117379 11661
rect 119200 11658 120000 11688
rect 117313 11656 120000 11658
rect 117313 11600 117318 11656
rect 117374 11600 120000 11656
rect 117313 11598 120000 11600
rect 117313 11595 117379 11598
rect 119200 11568 120000 11598
rect 15670 11456 15986 11457
rect 15670 11392 15676 11456
rect 15740 11392 15756 11456
rect 15820 11392 15836 11456
rect 15900 11392 15916 11456
rect 15980 11392 15986 11456
rect 15670 11391 15986 11392
rect 45118 11456 45434 11457
rect 45118 11392 45124 11456
rect 45188 11392 45204 11456
rect 45268 11392 45284 11456
rect 45348 11392 45364 11456
rect 45428 11392 45434 11456
rect 45118 11391 45434 11392
rect 74566 11456 74882 11457
rect 74566 11392 74572 11456
rect 74636 11392 74652 11456
rect 74716 11392 74732 11456
rect 74796 11392 74812 11456
rect 74876 11392 74882 11456
rect 74566 11391 74882 11392
rect 104014 11456 104330 11457
rect 104014 11392 104020 11456
rect 104084 11392 104100 11456
rect 104164 11392 104180 11456
rect 104244 11392 104260 11456
rect 104324 11392 104330 11456
rect 104014 11391 104330 11392
rect 117957 10978 118023 10981
rect 119200 10978 120000 11008
rect 117957 10976 120000 10978
rect 117957 10920 117962 10976
rect 118018 10920 120000 10976
rect 117957 10918 120000 10920
rect 117957 10915 118023 10918
rect 30394 10912 30710 10913
rect 30394 10848 30400 10912
rect 30464 10848 30480 10912
rect 30544 10848 30560 10912
rect 30624 10848 30640 10912
rect 30704 10848 30710 10912
rect 30394 10847 30710 10848
rect 59842 10912 60158 10913
rect 59842 10848 59848 10912
rect 59912 10848 59928 10912
rect 59992 10848 60008 10912
rect 60072 10848 60088 10912
rect 60152 10848 60158 10912
rect 59842 10847 60158 10848
rect 89290 10912 89606 10913
rect 89290 10848 89296 10912
rect 89360 10848 89376 10912
rect 89440 10848 89456 10912
rect 89520 10848 89536 10912
rect 89600 10848 89606 10912
rect 119200 10888 120000 10918
rect 89290 10847 89606 10848
rect 15670 10368 15986 10369
rect 0 10298 800 10328
rect 15670 10304 15676 10368
rect 15740 10304 15756 10368
rect 15820 10304 15836 10368
rect 15900 10304 15916 10368
rect 15980 10304 15986 10368
rect 15670 10303 15986 10304
rect 45118 10368 45434 10369
rect 45118 10304 45124 10368
rect 45188 10304 45204 10368
rect 45268 10304 45284 10368
rect 45348 10304 45364 10368
rect 45428 10304 45434 10368
rect 45118 10303 45434 10304
rect 74566 10368 74882 10369
rect 74566 10304 74572 10368
rect 74636 10304 74652 10368
rect 74716 10304 74732 10368
rect 74796 10304 74812 10368
rect 74876 10304 74882 10368
rect 74566 10303 74882 10304
rect 104014 10368 104330 10369
rect 104014 10304 104020 10368
rect 104084 10304 104100 10368
rect 104164 10304 104180 10368
rect 104244 10304 104260 10368
rect 104324 10304 104330 10368
rect 104014 10303 104330 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 30394 9824 30710 9825
rect 30394 9760 30400 9824
rect 30464 9760 30480 9824
rect 30544 9760 30560 9824
rect 30624 9760 30640 9824
rect 30704 9760 30710 9824
rect 30394 9759 30710 9760
rect 59842 9824 60158 9825
rect 59842 9760 59848 9824
rect 59912 9760 59928 9824
rect 59992 9760 60008 9824
rect 60072 9760 60088 9824
rect 60152 9760 60158 9824
rect 59842 9759 60158 9760
rect 89290 9824 89606 9825
rect 89290 9760 89296 9824
rect 89360 9760 89376 9824
rect 89440 9760 89456 9824
rect 89520 9760 89536 9824
rect 89600 9760 89606 9824
rect 89290 9759 89606 9760
rect 0 9618 800 9648
rect 1853 9618 1919 9621
rect 0 9616 1919 9618
rect 0 9560 1858 9616
rect 1914 9560 1919 9616
rect 0 9558 1919 9560
rect 0 9528 800 9558
rect 1853 9555 1919 9558
rect 117957 9618 118023 9621
rect 119200 9618 120000 9648
rect 117957 9616 120000 9618
rect 117957 9560 117962 9616
rect 118018 9560 120000 9616
rect 117957 9558 120000 9560
rect 117957 9555 118023 9558
rect 119200 9528 120000 9558
rect 15670 9280 15986 9281
rect 15670 9216 15676 9280
rect 15740 9216 15756 9280
rect 15820 9216 15836 9280
rect 15900 9216 15916 9280
rect 15980 9216 15986 9280
rect 15670 9215 15986 9216
rect 45118 9280 45434 9281
rect 45118 9216 45124 9280
rect 45188 9216 45204 9280
rect 45268 9216 45284 9280
rect 45348 9216 45364 9280
rect 45428 9216 45434 9280
rect 45118 9215 45434 9216
rect 74566 9280 74882 9281
rect 74566 9216 74572 9280
rect 74636 9216 74652 9280
rect 74716 9216 74732 9280
rect 74796 9216 74812 9280
rect 74876 9216 74882 9280
rect 74566 9215 74882 9216
rect 104014 9280 104330 9281
rect 104014 9216 104020 9280
rect 104084 9216 104100 9280
rect 104164 9216 104180 9280
rect 104244 9216 104260 9280
rect 104324 9216 104330 9280
rect 104014 9215 104330 9216
rect 115381 8938 115447 8941
rect 119200 8938 120000 8968
rect 115381 8936 120000 8938
rect 115381 8880 115386 8936
rect 115442 8880 120000 8936
rect 115381 8878 120000 8880
rect 115381 8875 115447 8878
rect 119200 8848 120000 8878
rect 30394 8736 30710 8737
rect 30394 8672 30400 8736
rect 30464 8672 30480 8736
rect 30544 8672 30560 8736
rect 30624 8672 30640 8736
rect 30704 8672 30710 8736
rect 30394 8671 30710 8672
rect 59842 8736 60158 8737
rect 59842 8672 59848 8736
rect 59912 8672 59928 8736
rect 59992 8672 60008 8736
rect 60072 8672 60088 8736
rect 60152 8672 60158 8736
rect 59842 8671 60158 8672
rect 89290 8736 89606 8737
rect 89290 8672 89296 8736
rect 89360 8672 89376 8736
rect 89440 8672 89456 8736
rect 89520 8672 89536 8736
rect 89600 8672 89606 8736
rect 89290 8671 89606 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 117957 8258 118023 8261
rect 119200 8258 120000 8288
rect 117957 8256 120000 8258
rect 117957 8200 117962 8256
rect 118018 8200 120000 8256
rect 117957 8198 120000 8200
rect 117957 8195 118023 8198
rect 15670 8192 15986 8193
rect 15670 8128 15676 8192
rect 15740 8128 15756 8192
rect 15820 8128 15836 8192
rect 15900 8128 15916 8192
rect 15980 8128 15986 8192
rect 15670 8127 15986 8128
rect 45118 8192 45434 8193
rect 45118 8128 45124 8192
rect 45188 8128 45204 8192
rect 45268 8128 45284 8192
rect 45348 8128 45364 8192
rect 45428 8128 45434 8192
rect 45118 8127 45434 8128
rect 74566 8192 74882 8193
rect 74566 8128 74572 8192
rect 74636 8128 74652 8192
rect 74716 8128 74732 8192
rect 74796 8128 74812 8192
rect 74876 8128 74882 8192
rect 74566 8127 74882 8128
rect 104014 8192 104330 8193
rect 104014 8128 104020 8192
rect 104084 8128 104100 8192
rect 104164 8128 104180 8192
rect 104244 8128 104260 8192
rect 104324 8128 104330 8192
rect 119200 8168 120000 8198
rect 104014 8127 104330 8128
rect 30394 7648 30710 7649
rect 0 7578 800 7608
rect 30394 7584 30400 7648
rect 30464 7584 30480 7648
rect 30544 7584 30560 7648
rect 30624 7584 30640 7648
rect 30704 7584 30710 7648
rect 30394 7583 30710 7584
rect 59842 7648 60158 7649
rect 59842 7584 59848 7648
rect 59912 7584 59928 7648
rect 59992 7584 60008 7648
rect 60072 7584 60088 7648
rect 60152 7584 60158 7648
rect 59842 7583 60158 7584
rect 89290 7648 89606 7649
rect 89290 7584 89296 7648
rect 89360 7584 89376 7648
rect 89440 7584 89456 7648
rect 89520 7584 89536 7648
rect 89600 7584 89606 7648
rect 89290 7583 89606 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 800 7518
rect 1393 7515 1459 7518
rect 15670 7104 15986 7105
rect 15670 7040 15676 7104
rect 15740 7040 15756 7104
rect 15820 7040 15836 7104
rect 15900 7040 15916 7104
rect 15980 7040 15986 7104
rect 15670 7039 15986 7040
rect 45118 7104 45434 7105
rect 45118 7040 45124 7104
rect 45188 7040 45204 7104
rect 45268 7040 45284 7104
rect 45348 7040 45364 7104
rect 45428 7040 45434 7104
rect 45118 7039 45434 7040
rect 74566 7104 74882 7105
rect 74566 7040 74572 7104
rect 74636 7040 74652 7104
rect 74716 7040 74732 7104
rect 74796 7040 74812 7104
rect 74876 7040 74882 7104
rect 74566 7039 74882 7040
rect 104014 7104 104330 7105
rect 104014 7040 104020 7104
rect 104084 7040 104100 7104
rect 104164 7040 104180 7104
rect 104244 7040 104260 7104
rect 104324 7040 104330 7104
rect 104014 7039 104330 7040
rect 117957 6898 118023 6901
rect 119200 6898 120000 6928
rect 117957 6896 120000 6898
rect 117957 6840 117962 6896
rect 118018 6840 120000 6896
rect 117957 6838 120000 6840
rect 117957 6835 118023 6838
rect 119200 6808 120000 6838
rect 30394 6560 30710 6561
rect 30394 6496 30400 6560
rect 30464 6496 30480 6560
rect 30544 6496 30560 6560
rect 30624 6496 30640 6560
rect 30704 6496 30710 6560
rect 30394 6495 30710 6496
rect 59842 6560 60158 6561
rect 59842 6496 59848 6560
rect 59912 6496 59928 6560
rect 59992 6496 60008 6560
rect 60072 6496 60088 6560
rect 60152 6496 60158 6560
rect 59842 6495 60158 6496
rect 89290 6560 89606 6561
rect 89290 6496 89296 6560
rect 89360 6496 89376 6560
rect 89440 6496 89456 6560
rect 89520 6496 89536 6560
rect 89600 6496 89606 6560
rect 89290 6495 89606 6496
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 117865 6218 117931 6221
rect 119200 6218 120000 6248
rect 117865 6216 120000 6218
rect 117865 6160 117870 6216
rect 117926 6160 120000 6216
rect 117865 6158 120000 6160
rect 117865 6155 117931 6158
rect 119200 6128 120000 6158
rect 15670 6016 15986 6017
rect 15670 5952 15676 6016
rect 15740 5952 15756 6016
rect 15820 5952 15836 6016
rect 15900 5952 15916 6016
rect 15980 5952 15986 6016
rect 15670 5951 15986 5952
rect 45118 6016 45434 6017
rect 45118 5952 45124 6016
rect 45188 5952 45204 6016
rect 45268 5952 45284 6016
rect 45348 5952 45364 6016
rect 45428 5952 45434 6016
rect 45118 5951 45434 5952
rect 74566 6016 74882 6017
rect 74566 5952 74572 6016
rect 74636 5952 74652 6016
rect 74716 5952 74732 6016
rect 74796 5952 74812 6016
rect 74876 5952 74882 6016
rect 74566 5951 74882 5952
rect 104014 6016 104330 6017
rect 104014 5952 104020 6016
rect 104084 5952 104100 6016
rect 104164 5952 104180 6016
rect 104244 5952 104260 6016
rect 104324 5952 104330 6016
rect 104014 5951 104330 5952
rect 0 5538 800 5568
rect 1853 5538 1919 5541
rect 0 5536 1919 5538
rect 0 5480 1858 5536
rect 1914 5480 1919 5536
rect 0 5478 1919 5480
rect 0 5448 800 5478
rect 1853 5475 1919 5478
rect 30394 5472 30710 5473
rect 30394 5408 30400 5472
rect 30464 5408 30480 5472
rect 30544 5408 30560 5472
rect 30624 5408 30640 5472
rect 30704 5408 30710 5472
rect 30394 5407 30710 5408
rect 59842 5472 60158 5473
rect 59842 5408 59848 5472
rect 59912 5408 59928 5472
rect 59992 5408 60008 5472
rect 60072 5408 60088 5472
rect 60152 5408 60158 5472
rect 59842 5407 60158 5408
rect 89290 5472 89606 5473
rect 89290 5408 89296 5472
rect 89360 5408 89376 5472
rect 89440 5408 89456 5472
rect 89520 5408 89536 5472
rect 89600 5408 89606 5472
rect 89290 5407 89606 5408
rect 15670 4928 15986 4929
rect 0 4858 800 4888
rect 15670 4864 15676 4928
rect 15740 4864 15756 4928
rect 15820 4864 15836 4928
rect 15900 4864 15916 4928
rect 15980 4864 15986 4928
rect 15670 4863 15986 4864
rect 45118 4928 45434 4929
rect 45118 4864 45124 4928
rect 45188 4864 45204 4928
rect 45268 4864 45284 4928
rect 45348 4864 45364 4928
rect 45428 4864 45434 4928
rect 45118 4863 45434 4864
rect 74566 4928 74882 4929
rect 74566 4864 74572 4928
rect 74636 4864 74652 4928
rect 74716 4864 74732 4928
rect 74796 4864 74812 4928
rect 74876 4864 74882 4928
rect 74566 4863 74882 4864
rect 104014 4928 104330 4929
rect 104014 4864 104020 4928
rect 104084 4864 104100 4928
rect 104164 4864 104180 4928
rect 104244 4864 104260 4928
rect 104324 4864 104330 4928
rect 104014 4863 104330 4864
rect 1393 4858 1459 4861
rect 0 4856 1459 4858
rect 0 4800 1398 4856
rect 1454 4800 1459 4856
rect 0 4798 1459 4800
rect 0 4768 800 4798
rect 1393 4795 1459 4798
rect 117957 4858 118023 4861
rect 119200 4858 120000 4888
rect 117957 4856 120000 4858
rect 117957 4800 117962 4856
rect 118018 4800 120000 4856
rect 117957 4798 120000 4800
rect 117957 4795 118023 4798
rect 119200 4768 120000 4798
rect 30394 4384 30710 4385
rect 30394 4320 30400 4384
rect 30464 4320 30480 4384
rect 30544 4320 30560 4384
rect 30624 4320 30640 4384
rect 30704 4320 30710 4384
rect 30394 4319 30710 4320
rect 59842 4384 60158 4385
rect 59842 4320 59848 4384
rect 59912 4320 59928 4384
rect 59992 4320 60008 4384
rect 60072 4320 60088 4384
rect 60152 4320 60158 4384
rect 59842 4319 60158 4320
rect 89290 4384 89606 4385
rect 89290 4320 89296 4384
rect 89360 4320 89376 4384
rect 89440 4320 89456 4384
rect 89520 4320 89536 4384
rect 89600 4320 89606 4384
rect 89290 4319 89606 4320
rect 117773 4178 117839 4181
rect 119200 4178 120000 4208
rect 117773 4176 120000 4178
rect 117773 4120 117778 4176
rect 117834 4120 120000 4176
rect 117773 4118 120000 4120
rect 117773 4115 117839 4118
rect 119200 4088 120000 4118
rect 15670 3840 15986 3841
rect 15670 3776 15676 3840
rect 15740 3776 15756 3840
rect 15820 3776 15836 3840
rect 15900 3776 15916 3840
rect 15980 3776 15986 3840
rect 15670 3775 15986 3776
rect 45118 3840 45434 3841
rect 45118 3776 45124 3840
rect 45188 3776 45204 3840
rect 45268 3776 45284 3840
rect 45348 3776 45364 3840
rect 45428 3776 45434 3840
rect 45118 3775 45434 3776
rect 74566 3840 74882 3841
rect 74566 3776 74572 3840
rect 74636 3776 74652 3840
rect 74716 3776 74732 3840
rect 74796 3776 74812 3840
rect 74876 3776 74882 3840
rect 74566 3775 74882 3776
rect 104014 3840 104330 3841
rect 104014 3776 104020 3840
rect 104084 3776 104100 3840
rect 104164 3776 104180 3840
rect 104244 3776 104260 3840
rect 104324 3776 104330 3840
rect 104014 3775 104330 3776
rect 57973 3770 58039 3773
rect 59629 3770 59695 3773
rect 57973 3768 59695 3770
rect 57973 3712 57978 3768
rect 58034 3712 59634 3768
rect 59690 3712 59695 3768
rect 57973 3710 59695 3712
rect 57973 3707 58039 3710
rect 59629 3707 59695 3710
rect 40309 3634 40375 3637
rect 47301 3634 47367 3637
rect 40309 3632 47367 3634
rect 40309 3576 40314 3632
rect 40370 3576 47306 3632
rect 47362 3576 47367 3632
rect 40309 3574 47367 3576
rect 40309 3571 40375 3574
rect 47301 3571 47367 3574
rect 58065 3634 58131 3637
rect 58525 3634 58591 3637
rect 58065 3632 58591 3634
rect 58065 3576 58070 3632
rect 58126 3576 58530 3632
rect 58586 3576 58591 3632
rect 58065 3574 58591 3576
rect 58065 3571 58131 3574
rect 58525 3571 58591 3574
rect 0 3498 800 3528
rect 1577 3498 1643 3501
rect 0 3496 1643 3498
rect 0 3440 1582 3496
rect 1638 3440 1643 3496
rect 0 3438 1643 3440
rect 0 3408 800 3438
rect 1577 3435 1643 3438
rect 42425 3498 42491 3501
rect 48037 3498 48103 3501
rect 42425 3496 48103 3498
rect 42425 3440 42430 3496
rect 42486 3440 48042 3496
rect 48098 3440 48103 3496
rect 42425 3438 48103 3440
rect 42425 3435 42491 3438
rect 48037 3435 48103 3438
rect 43253 3362 43319 3365
rect 47577 3362 47643 3365
rect 43253 3360 47643 3362
rect 43253 3304 43258 3360
rect 43314 3304 47582 3360
rect 47638 3304 47643 3360
rect 43253 3302 47643 3304
rect 43253 3299 43319 3302
rect 47577 3299 47643 3302
rect 30394 3296 30710 3297
rect 30394 3232 30400 3296
rect 30464 3232 30480 3296
rect 30544 3232 30560 3296
rect 30624 3232 30640 3296
rect 30704 3232 30710 3296
rect 30394 3231 30710 3232
rect 59842 3296 60158 3297
rect 59842 3232 59848 3296
rect 59912 3232 59928 3296
rect 59992 3232 60008 3296
rect 60072 3232 60088 3296
rect 60152 3232 60158 3296
rect 59842 3231 60158 3232
rect 89290 3296 89606 3297
rect 89290 3232 89296 3296
rect 89360 3232 89376 3296
rect 89440 3232 89456 3296
rect 89520 3232 89536 3296
rect 89600 3232 89606 3296
rect 89290 3231 89606 3232
rect 41229 3226 41295 3229
rect 46197 3226 46263 3229
rect 41229 3224 46263 3226
rect 41229 3168 41234 3224
rect 41290 3168 46202 3224
rect 46258 3168 46263 3224
rect 41229 3166 46263 3168
rect 41229 3163 41295 3166
rect 46197 3163 46263 3166
rect 57237 3226 57303 3229
rect 58065 3226 58131 3229
rect 57237 3224 58131 3226
rect 57237 3168 57242 3224
rect 57298 3168 58070 3224
rect 58126 3168 58131 3224
rect 57237 3166 58131 3168
rect 57237 3163 57303 3166
rect 58065 3163 58131 3166
rect 40033 3090 40099 3093
rect 45369 3090 45435 3093
rect 40033 3088 45435 3090
rect 40033 3032 40038 3088
rect 40094 3032 45374 3088
rect 45430 3032 45435 3088
rect 40033 3030 45435 3032
rect 40033 3027 40099 3030
rect 45369 3027 45435 3030
rect 57697 3090 57763 3093
rect 66161 3090 66227 3093
rect 57697 3088 66227 3090
rect 57697 3032 57702 3088
rect 57758 3032 66166 3088
rect 66222 3032 66227 3088
rect 57697 3030 66227 3032
rect 57697 3027 57763 3030
rect 66161 3027 66227 3030
rect 70301 3090 70367 3093
rect 77109 3090 77175 3093
rect 70301 3088 77175 3090
rect 70301 3032 70306 3088
rect 70362 3032 77114 3088
rect 77170 3032 77175 3088
rect 70301 3030 77175 3032
rect 70301 3027 70367 3030
rect 77109 3027 77175 3030
rect 39849 2954 39915 2957
rect 47485 2954 47551 2957
rect 39849 2952 47551 2954
rect 39849 2896 39854 2952
rect 39910 2896 47490 2952
rect 47546 2896 47551 2952
rect 39849 2894 47551 2896
rect 39849 2891 39915 2894
rect 47485 2891 47551 2894
rect 55581 2954 55647 2957
rect 57789 2954 57855 2957
rect 55581 2952 57855 2954
rect 55581 2896 55586 2952
rect 55642 2896 57794 2952
rect 57850 2896 57855 2952
rect 55581 2894 57855 2896
rect 55581 2891 55647 2894
rect 57789 2891 57855 2894
rect 58709 2954 58775 2957
rect 64045 2954 64111 2957
rect 58709 2952 64111 2954
rect 58709 2896 58714 2952
rect 58770 2896 64050 2952
rect 64106 2896 64111 2952
rect 58709 2894 64111 2896
rect 58709 2891 58775 2894
rect 64045 2891 64111 2894
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 57973 2818 58039 2821
rect 58801 2818 58867 2821
rect 57973 2816 58867 2818
rect 57973 2760 57978 2816
rect 58034 2760 58806 2816
rect 58862 2760 58867 2816
rect 57973 2758 58867 2760
rect 57973 2755 58039 2758
rect 58801 2755 58867 2758
rect 60917 2818 60983 2821
rect 73429 2818 73495 2821
rect 60917 2816 73495 2818
rect 60917 2760 60922 2816
rect 60978 2760 73434 2816
rect 73490 2760 73495 2816
rect 60917 2758 73495 2760
rect 60917 2755 60983 2758
rect 73429 2755 73495 2758
rect 77201 2818 77267 2821
rect 78029 2818 78095 2821
rect 77201 2816 78095 2818
rect 77201 2760 77206 2816
rect 77262 2760 78034 2816
rect 78090 2760 78095 2816
rect 77201 2758 78095 2760
rect 77201 2755 77267 2758
rect 78029 2755 78095 2758
rect 117865 2818 117931 2821
rect 119200 2818 120000 2848
rect 117865 2816 120000 2818
rect 117865 2760 117870 2816
rect 117926 2760 120000 2816
rect 117865 2758 120000 2760
rect 117865 2755 117931 2758
rect 15670 2752 15986 2753
rect 15670 2688 15676 2752
rect 15740 2688 15756 2752
rect 15820 2688 15836 2752
rect 15900 2688 15916 2752
rect 15980 2688 15986 2752
rect 15670 2687 15986 2688
rect 45118 2752 45434 2753
rect 45118 2688 45124 2752
rect 45188 2688 45204 2752
rect 45268 2688 45284 2752
rect 45348 2688 45364 2752
rect 45428 2688 45434 2752
rect 45118 2687 45434 2688
rect 74566 2752 74882 2753
rect 74566 2688 74572 2752
rect 74636 2688 74652 2752
rect 74716 2688 74732 2752
rect 74796 2688 74812 2752
rect 74876 2688 74882 2752
rect 74566 2687 74882 2688
rect 104014 2752 104330 2753
rect 104014 2688 104020 2752
rect 104084 2688 104100 2752
rect 104164 2688 104180 2752
rect 104244 2688 104260 2752
rect 104324 2688 104330 2752
rect 119200 2728 120000 2758
rect 104014 2687 104330 2688
rect 55489 2682 55555 2685
rect 62573 2682 62639 2685
rect 55489 2680 62639 2682
rect 55489 2624 55494 2680
rect 55550 2624 62578 2680
rect 62634 2624 62639 2680
rect 55489 2622 62639 2624
rect 55489 2619 55555 2622
rect 62573 2619 62639 2622
rect 62757 2682 62823 2685
rect 67265 2682 67331 2685
rect 62757 2680 67331 2682
rect 62757 2624 62762 2680
rect 62818 2624 67270 2680
rect 67326 2624 67331 2680
rect 62757 2622 67331 2624
rect 62757 2619 62823 2622
rect 67265 2619 67331 2622
rect 16849 2546 16915 2549
rect 74625 2546 74691 2549
rect 16849 2544 74691 2546
rect 16849 2488 16854 2544
rect 16910 2488 74630 2544
rect 74686 2488 74691 2544
rect 16849 2486 74691 2488
rect 16849 2483 16915 2486
rect 74625 2483 74691 2486
rect 89529 2546 89595 2549
rect 92197 2546 92263 2549
rect 89529 2544 92263 2546
rect 89529 2488 89534 2544
rect 89590 2488 92202 2544
rect 92258 2488 92263 2544
rect 89529 2486 92263 2488
rect 89529 2483 89595 2486
rect 92197 2483 92263 2486
rect 19701 2410 19767 2413
rect 28165 2410 28231 2413
rect 19701 2408 28231 2410
rect 19701 2352 19706 2408
rect 19762 2352 28170 2408
rect 28226 2352 28231 2408
rect 19701 2350 28231 2352
rect 19701 2347 19767 2350
rect 28165 2347 28231 2350
rect 39573 2410 39639 2413
rect 46749 2410 46815 2413
rect 39573 2408 46815 2410
rect 39573 2352 39578 2408
rect 39634 2352 46754 2408
rect 46810 2352 46815 2408
rect 39573 2350 46815 2352
rect 39573 2347 39639 2350
rect 46749 2347 46815 2350
rect 47945 2410 48011 2413
rect 115565 2410 115631 2413
rect 47945 2408 115631 2410
rect 47945 2352 47950 2408
rect 48006 2352 115570 2408
rect 115626 2352 115631 2408
rect 47945 2350 115631 2352
rect 47945 2347 48011 2350
rect 115565 2347 115631 2350
rect 61009 2274 61075 2277
rect 69933 2274 69999 2277
rect 61009 2272 69999 2274
rect 61009 2216 61014 2272
rect 61070 2216 69938 2272
rect 69994 2216 69999 2272
rect 61009 2214 69999 2216
rect 61009 2211 61075 2214
rect 69933 2211 69999 2214
rect 70669 2274 70735 2277
rect 79593 2274 79659 2277
rect 80145 2274 80211 2277
rect 70669 2272 77310 2274
rect 70669 2216 70674 2272
rect 70730 2216 77310 2272
rect 70669 2214 77310 2216
rect 70669 2211 70735 2214
rect 30394 2208 30710 2209
rect 30394 2144 30400 2208
rect 30464 2144 30480 2208
rect 30544 2144 30560 2208
rect 30624 2144 30640 2208
rect 30704 2144 30710 2208
rect 30394 2143 30710 2144
rect 59842 2208 60158 2209
rect 59842 2144 59848 2208
rect 59912 2144 59928 2208
rect 59992 2144 60008 2208
rect 60072 2144 60088 2208
rect 60152 2144 60158 2208
rect 59842 2143 60158 2144
rect 51993 2138 52059 2141
rect 53833 2138 53899 2141
rect 55305 2138 55371 2141
rect 51993 2136 55371 2138
rect 51993 2080 51998 2136
rect 52054 2080 53838 2136
rect 53894 2080 55310 2136
rect 55366 2080 55371 2136
rect 51993 2078 55371 2080
rect 51993 2075 52059 2078
rect 53833 2075 53899 2078
rect 55305 2075 55371 2078
rect 60641 2138 60707 2141
rect 67449 2138 67515 2141
rect 60641 2136 67515 2138
rect 60641 2080 60646 2136
rect 60702 2080 67454 2136
rect 67510 2080 67515 2136
rect 60641 2078 67515 2080
rect 77250 2138 77310 2214
rect 79593 2272 80211 2274
rect 79593 2216 79598 2272
rect 79654 2216 80150 2272
rect 80206 2216 80211 2272
rect 79593 2214 80211 2216
rect 79593 2211 79659 2214
rect 80145 2211 80211 2214
rect 89290 2208 89606 2209
rect 89290 2144 89296 2208
rect 89360 2144 89376 2208
rect 89440 2144 89456 2208
rect 89520 2144 89536 2208
rect 89600 2144 89606 2208
rect 89290 2143 89606 2144
rect 89713 2138 89779 2141
rect 92289 2138 92355 2141
rect 77250 2078 86970 2138
rect 60641 2075 60707 2078
rect 67449 2075 67515 2078
rect 55213 2002 55279 2005
rect 61009 2002 61075 2005
rect 55213 2000 61075 2002
rect 55213 1944 55218 2000
rect 55274 1944 61014 2000
rect 61070 1944 61075 2000
rect 55213 1942 61075 1944
rect 55213 1939 55279 1942
rect 61009 1939 61075 1942
rect 72325 2002 72391 2005
rect 77385 2002 77451 2005
rect 72325 2000 77451 2002
rect 72325 1944 72330 2000
rect 72386 1944 77390 2000
rect 77446 1944 77451 2000
rect 72325 1942 77451 1944
rect 72325 1939 72391 1942
rect 77385 1939 77451 1942
rect 30741 1866 30807 1869
rect 38561 1866 38627 1869
rect 30741 1864 38627 1866
rect 30741 1808 30746 1864
rect 30802 1808 38566 1864
rect 38622 1808 38627 1864
rect 30741 1806 38627 1808
rect 30741 1803 30807 1806
rect 38561 1803 38627 1806
rect 58157 1866 58223 1869
rect 67357 1866 67423 1869
rect 58157 1864 67423 1866
rect 58157 1808 58162 1864
rect 58218 1808 67362 1864
rect 67418 1808 67423 1864
rect 58157 1806 67423 1808
rect 58157 1803 58223 1806
rect 67357 1803 67423 1806
rect 70945 1866 71011 1869
rect 75545 1866 75611 1869
rect 70945 1864 75611 1866
rect 70945 1808 70950 1864
rect 71006 1808 75550 1864
rect 75606 1808 75611 1864
rect 70945 1806 75611 1808
rect 70945 1803 71011 1806
rect 75545 1803 75611 1806
rect 26141 1730 26207 1733
rect 31569 1730 31635 1733
rect 26141 1728 31635 1730
rect 26141 1672 26146 1728
rect 26202 1672 31574 1728
rect 31630 1672 31635 1728
rect 26141 1670 31635 1672
rect 26141 1667 26207 1670
rect 31569 1667 31635 1670
rect 58065 1730 58131 1733
rect 60825 1730 60891 1733
rect 58065 1728 60891 1730
rect 58065 1672 58070 1728
rect 58126 1672 60830 1728
rect 60886 1672 60891 1728
rect 58065 1670 60891 1672
rect 58065 1667 58131 1670
rect 60825 1667 60891 1670
rect 61285 1730 61351 1733
rect 64137 1730 64203 1733
rect 66897 1730 66963 1733
rect 61285 1728 66963 1730
rect 61285 1672 61290 1728
rect 61346 1672 64142 1728
rect 64198 1672 66902 1728
rect 66958 1672 66963 1728
rect 61285 1670 66963 1672
rect 61285 1667 61351 1670
rect 64137 1667 64203 1670
rect 66897 1667 66963 1670
rect 72877 1730 72943 1733
rect 77845 1730 77911 1733
rect 72877 1728 77911 1730
rect 72877 1672 72882 1728
rect 72938 1672 77850 1728
rect 77906 1672 77911 1728
rect 72877 1670 77911 1672
rect 86910 1730 86970 2078
rect 89713 2136 92355 2138
rect 89713 2080 89718 2136
rect 89774 2080 92294 2136
rect 92350 2080 92355 2136
rect 89713 2078 92355 2080
rect 89713 2075 89779 2078
rect 92289 2075 92355 2078
rect 116393 2138 116459 2141
rect 119200 2138 120000 2168
rect 116393 2136 120000 2138
rect 116393 2080 116398 2136
rect 116454 2080 120000 2136
rect 116393 2078 120000 2080
rect 116393 2075 116459 2078
rect 119200 2048 120000 2078
rect 89437 1866 89503 1869
rect 89805 1866 89871 1869
rect 89437 1864 89871 1866
rect 89437 1808 89442 1864
rect 89498 1808 89810 1864
rect 89866 1808 89871 1864
rect 89437 1806 89871 1808
rect 89437 1803 89503 1806
rect 89805 1803 89871 1806
rect 89621 1730 89687 1733
rect 86910 1728 89687 1730
rect 86910 1672 89626 1728
rect 89682 1672 89687 1728
rect 86910 1670 89687 1672
rect 72877 1667 72943 1670
rect 77845 1667 77911 1670
rect 89621 1667 89687 1670
rect 17309 1594 17375 1597
rect 28441 1594 28507 1597
rect 17309 1592 28507 1594
rect 17309 1536 17314 1592
rect 17370 1536 28446 1592
rect 28502 1536 28507 1592
rect 17309 1534 28507 1536
rect 17309 1531 17375 1534
rect 28441 1531 28507 1534
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 80053 1458 80119 1461
rect 88977 1458 89043 1461
rect 80053 1456 89043 1458
rect 80053 1400 80058 1456
rect 80114 1400 88982 1456
rect 89038 1400 89043 1456
rect 80053 1398 89043 1400
rect 80053 1395 80119 1398
rect 88977 1395 89043 1398
rect 89345 1458 89411 1461
rect 90909 1458 90975 1461
rect 89345 1456 90975 1458
rect 89345 1400 89350 1456
rect 89406 1400 90914 1456
rect 90970 1400 90975 1456
rect 89345 1398 90975 1400
rect 89345 1395 89411 1398
rect 90909 1395 90975 1398
rect 116669 1458 116735 1461
rect 119200 1458 120000 1488
rect 116669 1456 120000 1458
rect 116669 1400 116674 1456
rect 116730 1400 120000 1456
rect 116669 1398 120000 1400
rect 116669 1395 116735 1398
rect 119200 1368 120000 1398
rect 0 778 800 808
rect 1393 778 1459 781
rect 0 776 1459 778
rect 0 720 1398 776
rect 1454 720 1459 776
rect 0 718 1459 720
rect 0 688 800 718
rect 1393 715 1459 718
rect 117773 98 117839 101
rect 119200 98 120000 128
rect 117773 96 120000 98
rect 117773 40 117778 96
rect 117834 40 120000 96
rect 117773 38 120000 40
rect 117773 35 117839 38
rect 119200 8 120000 38
<< via3 >>
rect 15676 27772 15740 27776
rect 15676 27716 15680 27772
rect 15680 27716 15736 27772
rect 15736 27716 15740 27772
rect 15676 27712 15740 27716
rect 15756 27772 15820 27776
rect 15756 27716 15760 27772
rect 15760 27716 15816 27772
rect 15816 27716 15820 27772
rect 15756 27712 15820 27716
rect 15836 27772 15900 27776
rect 15836 27716 15840 27772
rect 15840 27716 15896 27772
rect 15896 27716 15900 27772
rect 15836 27712 15900 27716
rect 15916 27772 15980 27776
rect 15916 27716 15920 27772
rect 15920 27716 15976 27772
rect 15976 27716 15980 27772
rect 15916 27712 15980 27716
rect 45124 27772 45188 27776
rect 45124 27716 45128 27772
rect 45128 27716 45184 27772
rect 45184 27716 45188 27772
rect 45124 27712 45188 27716
rect 45204 27772 45268 27776
rect 45204 27716 45208 27772
rect 45208 27716 45264 27772
rect 45264 27716 45268 27772
rect 45204 27712 45268 27716
rect 45284 27772 45348 27776
rect 45284 27716 45288 27772
rect 45288 27716 45344 27772
rect 45344 27716 45348 27772
rect 45284 27712 45348 27716
rect 45364 27772 45428 27776
rect 45364 27716 45368 27772
rect 45368 27716 45424 27772
rect 45424 27716 45428 27772
rect 45364 27712 45428 27716
rect 74572 27772 74636 27776
rect 74572 27716 74576 27772
rect 74576 27716 74632 27772
rect 74632 27716 74636 27772
rect 74572 27712 74636 27716
rect 74652 27772 74716 27776
rect 74652 27716 74656 27772
rect 74656 27716 74712 27772
rect 74712 27716 74716 27772
rect 74652 27712 74716 27716
rect 74732 27772 74796 27776
rect 74732 27716 74736 27772
rect 74736 27716 74792 27772
rect 74792 27716 74796 27772
rect 74732 27712 74796 27716
rect 74812 27772 74876 27776
rect 74812 27716 74816 27772
rect 74816 27716 74872 27772
rect 74872 27716 74876 27772
rect 74812 27712 74876 27716
rect 104020 27772 104084 27776
rect 104020 27716 104024 27772
rect 104024 27716 104080 27772
rect 104080 27716 104084 27772
rect 104020 27712 104084 27716
rect 104100 27772 104164 27776
rect 104100 27716 104104 27772
rect 104104 27716 104160 27772
rect 104160 27716 104164 27772
rect 104100 27712 104164 27716
rect 104180 27772 104244 27776
rect 104180 27716 104184 27772
rect 104184 27716 104240 27772
rect 104240 27716 104244 27772
rect 104180 27712 104244 27716
rect 104260 27772 104324 27776
rect 104260 27716 104264 27772
rect 104264 27716 104320 27772
rect 104320 27716 104324 27772
rect 104260 27712 104324 27716
rect 30400 27228 30464 27232
rect 30400 27172 30404 27228
rect 30404 27172 30460 27228
rect 30460 27172 30464 27228
rect 30400 27168 30464 27172
rect 30480 27228 30544 27232
rect 30480 27172 30484 27228
rect 30484 27172 30540 27228
rect 30540 27172 30544 27228
rect 30480 27168 30544 27172
rect 30560 27228 30624 27232
rect 30560 27172 30564 27228
rect 30564 27172 30620 27228
rect 30620 27172 30624 27228
rect 30560 27168 30624 27172
rect 30640 27228 30704 27232
rect 30640 27172 30644 27228
rect 30644 27172 30700 27228
rect 30700 27172 30704 27228
rect 30640 27168 30704 27172
rect 59848 27228 59912 27232
rect 59848 27172 59852 27228
rect 59852 27172 59908 27228
rect 59908 27172 59912 27228
rect 59848 27168 59912 27172
rect 59928 27228 59992 27232
rect 59928 27172 59932 27228
rect 59932 27172 59988 27228
rect 59988 27172 59992 27228
rect 59928 27168 59992 27172
rect 60008 27228 60072 27232
rect 60008 27172 60012 27228
rect 60012 27172 60068 27228
rect 60068 27172 60072 27228
rect 60008 27168 60072 27172
rect 60088 27228 60152 27232
rect 60088 27172 60092 27228
rect 60092 27172 60148 27228
rect 60148 27172 60152 27228
rect 60088 27168 60152 27172
rect 89296 27228 89360 27232
rect 89296 27172 89300 27228
rect 89300 27172 89356 27228
rect 89356 27172 89360 27228
rect 89296 27168 89360 27172
rect 89376 27228 89440 27232
rect 89376 27172 89380 27228
rect 89380 27172 89436 27228
rect 89436 27172 89440 27228
rect 89376 27168 89440 27172
rect 89456 27228 89520 27232
rect 89456 27172 89460 27228
rect 89460 27172 89516 27228
rect 89516 27172 89520 27228
rect 89456 27168 89520 27172
rect 89536 27228 89600 27232
rect 89536 27172 89540 27228
rect 89540 27172 89596 27228
rect 89596 27172 89600 27228
rect 89536 27168 89600 27172
rect 70348 26692 70412 26756
rect 15676 26684 15740 26688
rect 15676 26628 15680 26684
rect 15680 26628 15736 26684
rect 15736 26628 15740 26684
rect 15676 26624 15740 26628
rect 15756 26684 15820 26688
rect 15756 26628 15760 26684
rect 15760 26628 15816 26684
rect 15816 26628 15820 26684
rect 15756 26624 15820 26628
rect 15836 26684 15900 26688
rect 15836 26628 15840 26684
rect 15840 26628 15896 26684
rect 15896 26628 15900 26684
rect 15836 26624 15900 26628
rect 15916 26684 15980 26688
rect 15916 26628 15920 26684
rect 15920 26628 15976 26684
rect 15976 26628 15980 26684
rect 15916 26624 15980 26628
rect 45124 26684 45188 26688
rect 45124 26628 45128 26684
rect 45128 26628 45184 26684
rect 45184 26628 45188 26684
rect 45124 26624 45188 26628
rect 45204 26684 45268 26688
rect 45204 26628 45208 26684
rect 45208 26628 45264 26684
rect 45264 26628 45268 26684
rect 45204 26624 45268 26628
rect 45284 26684 45348 26688
rect 45284 26628 45288 26684
rect 45288 26628 45344 26684
rect 45344 26628 45348 26684
rect 45284 26624 45348 26628
rect 45364 26684 45428 26688
rect 45364 26628 45368 26684
rect 45368 26628 45424 26684
rect 45424 26628 45428 26684
rect 45364 26624 45428 26628
rect 74572 26684 74636 26688
rect 74572 26628 74576 26684
rect 74576 26628 74632 26684
rect 74632 26628 74636 26684
rect 74572 26624 74636 26628
rect 74652 26684 74716 26688
rect 74652 26628 74656 26684
rect 74656 26628 74712 26684
rect 74712 26628 74716 26684
rect 74652 26624 74716 26628
rect 74732 26684 74796 26688
rect 74732 26628 74736 26684
rect 74736 26628 74792 26684
rect 74792 26628 74796 26684
rect 74732 26624 74796 26628
rect 74812 26684 74876 26688
rect 74812 26628 74816 26684
rect 74816 26628 74872 26684
rect 74872 26628 74876 26684
rect 74812 26624 74876 26628
rect 104020 26684 104084 26688
rect 104020 26628 104024 26684
rect 104024 26628 104080 26684
rect 104080 26628 104084 26684
rect 104020 26624 104084 26628
rect 104100 26684 104164 26688
rect 104100 26628 104104 26684
rect 104104 26628 104160 26684
rect 104160 26628 104164 26684
rect 104100 26624 104164 26628
rect 104180 26684 104244 26688
rect 104180 26628 104184 26684
rect 104184 26628 104240 26684
rect 104240 26628 104244 26684
rect 104180 26624 104244 26628
rect 104260 26684 104324 26688
rect 104260 26628 104264 26684
rect 104264 26628 104320 26684
rect 104320 26628 104324 26684
rect 104260 26624 104324 26628
rect 70716 26284 70780 26348
rect 30400 26140 30464 26144
rect 30400 26084 30404 26140
rect 30404 26084 30460 26140
rect 30460 26084 30464 26140
rect 30400 26080 30464 26084
rect 30480 26140 30544 26144
rect 30480 26084 30484 26140
rect 30484 26084 30540 26140
rect 30540 26084 30544 26140
rect 30480 26080 30544 26084
rect 30560 26140 30624 26144
rect 30560 26084 30564 26140
rect 30564 26084 30620 26140
rect 30620 26084 30624 26140
rect 30560 26080 30624 26084
rect 30640 26140 30704 26144
rect 30640 26084 30644 26140
rect 30644 26084 30700 26140
rect 30700 26084 30704 26140
rect 30640 26080 30704 26084
rect 59848 26140 59912 26144
rect 59848 26084 59852 26140
rect 59852 26084 59908 26140
rect 59908 26084 59912 26140
rect 59848 26080 59912 26084
rect 59928 26140 59992 26144
rect 59928 26084 59932 26140
rect 59932 26084 59988 26140
rect 59988 26084 59992 26140
rect 59928 26080 59992 26084
rect 60008 26140 60072 26144
rect 60008 26084 60012 26140
rect 60012 26084 60068 26140
rect 60068 26084 60072 26140
rect 60008 26080 60072 26084
rect 60088 26140 60152 26144
rect 60088 26084 60092 26140
rect 60092 26084 60148 26140
rect 60148 26084 60152 26140
rect 60088 26080 60152 26084
rect 89296 26140 89360 26144
rect 89296 26084 89300 26140
rect 89300 26084 89356 26140
rect 89356 26084 89360 26140
rect 89296 26080 89360 26084
rect 89376 26140 89440 26144
rect 89376 26084 89380 26140
rect 89380 26084 89436 26140
rect 89436 26084 89440 26140
rect 89376 26080 89440 26084
rect 89456 26140 89520 26144
rect 89456 26084 89460 26140
rect 89460 26084 89516 26140
rect 89516 26084 89520 26140
rect 89456 26080 89520 26084
rect 89536 26140 89600 26144
rect 89536 26084 89540 26140
rect 89540 26084 89596 26140
rect 89596 26084 89600 26140
rect 89536 26080 89600 26084
rect 15676 25596 15740 25600
rect 15676 25540 15680 25596
rect 15680 25540 15736 25596
rect 15736 25540 15740 25596
rect 15676 25536 15740 25540
rect 15756 25596 15820 25600
rect 15756 25540 15760 25596
rect 15760 25540 15816 25596
rect 15816 25540 15820 25596
rect 15756 25536 15820 25540
rect 15836 25596 15900 25600
rect 15836 25540 15840 25596
rect 15840 25540 15896 25596
rect 15896 25540 15900 25596
rect 15836 25536 15900 25540
rect 15916 25596 15980 25600
rect 15916 25540 15920 25596
rect 15920 25540 15976 25596
rect 15976 25540 15980 25596
rect 15916 25536 15980 25540
rect 45124 25596 45188 25600
rect 45124 25540 45128 25596
rect 45128 25540 45184 25596
rect 45184 25540 45188 25596
rect 45124 25536 45188 25540
rect 45204 25596 45268 25600
rect 45204 25540 45208 25596
rect 45208 25540 45264 25596
rect 45264 25540 45268 25596
rect 45204 25536 45268 25540
rect 45284 25596 45348 25600
rect 45284 25540 45288 25596
rect 45288 25540 45344 25596
rect 45344 25540 45348 25596
rect 45284 25536 45348 25540
rect 45364 25596 45428 25600
rect 45364 25540 45368 25596
rect 45368 25540 45424 25596
rect 45424 25540 45428 25596
rect 45364 25536 45428 25540
rect 74572 25596 74636 25600
rect 74572 25540 74576 25596
rect 74576 25540 74632 25596
rect 74632 25540 74636 25596
rect 74572 25536 74636 25540
rect 74652 25596 74716 25600
rect 74652 25540 74656 25596
rect 74656 25540 74712 25596
rect 74712 25540 74716 25596
rect 74652 25536 74716 25540
rect 74732 25596 74796 25600
rect 74732 25540 74736 25596
rect 74736 25540 74792 25596
rect 74792 25540 74796 25596
rect 74732 25536 74796 25540
rect 74812 25596 74876 25600
rect 74812 25540 74816 25596
rect 74816 25540 74872 25596
rect 74872 25540 74876 25596
rect 74812 25536 74876 25540
rect 104020 25596 104084 25600
rect 104020 25540 104024 25596
rect 104024 25540 104080 25596
rect 104080 25540 104084 25596
rect 104020 25536 104084 25540
rect 104100 25596 104164 25600
rect 104100 25540 104104 25596
rect 104104 25540 104160 25596
rect 104160 25540 104164 25596
rect 104100 25536 104164 25540
rect 104180 25596 104244 25600
rect 104180 25540 104184 25596
rect 104184 25540 104240 25596
rect 104240 25540 104244 25596
rect 104180 25536 104244 25540
rect 104260 25596 104324 25600
rect 104260 25540 104264 25596
rect 104264 25540 104320 25596
rect 104320 25540 104324 25596
rect 104260 25536 104324 25540
rect 30400 25052 30464 25056
rect 30400 24996 30404 25052
rect 30404 24996 30460 25052
rect 30460 24996 30464 25052
rect 30400 24992 30464 24996
rect 30480 25052 30544 25056
rect 30480 24996 30484 25052
rect 30484 24996 30540 25052
rect 30540 24996 30544 25052
rect 30480 24992 30544 24996
rect 30560 25052 30624 25056
rect 30560 24996 30564 25052
rect 30564 24996 30620 25052
rect 30620 24996 30624 25052
rect 30560 24992 30624 24996
rect 30640 25052 30704 25056
rect 30640 24996 30644 25052
rect 30644 24996 30700 25052
rect 30700 24996 30704 25052
rect 30640 24992 30704 24996
rect 59848 25052 59912 25056
rect 59848 24996 59852 25052
rect 59852 24996 59908 25052
rect 59908 24996 59912 25052
rect 59848 24992 59912 24996
rect 59928 25052 59992 25056
rect 59928 24996 59932 25052
rect 59932 24996 59988 25052
rect 59988 24996 59992 25052
rect 59928 24992 59992 24996
rect 60008 25052 60072 25056
rect 60008 24996 60012 25052
rect 60012 24996 60068 25052
rect 60068 24996 60072 25052
rect 60008 24992 60072 24996
rect 60088 25052 60152 25056
rect 60088 24996 60092 25052
rect 60092 24996 60148 25052
rect 60148 24996 60152 25052
rect 60088 24992 60152 24996
rect 89296 25052 89360 25056
rect 89296 24996 89300 25052
rect 89300 24996 89356 25052
rect 89356 24996 89360 25052
rect 89296 24992 89360 24996
rect 89376 25052 89440 25056
rect 89376 24996 89380 25052
rect 89380 24996 89436 25052
rect 89436 24996 89440 25052
rect 89376 24992 89440 24996
rect 89456 25052 89520 25056
rect 89456 24996 89460 25052
rect 89460 24996 89516 25052
rect 89516 24996 89520 25052
rect 89456 24992 89520 24996
rect 89536 25052 89600 25056
rect 89536 24996 89540 25052
rect 89540 24996 89596 25052
rect 89596 24996 89600 25052
rect 89536 24992 89600 24996
rect 15676 24508 15740 24512
rect 15676 24452 15680 24508
rect 15680 24452 15736 24508
rect 15736 24452 15740 24508
rect 15676 24448 15740 24452
rect 15756 24508 15820 24512
rect 15756 24452 15760 24508
rect 15760 24452 15816 24508
rect 15816 24452 15820 24508
rect 15756 24448 15820 24452
rect 15836 24508 15900 24512
rect 15836 24452 15840 24508
rect 15840 24452 15896 24508
rect 15896 24452 15900 24508
rect 15836 24448 15900 24452
rect 15916 24508 15980 24512
rect 15916 24452 15920 24508
rect 15920 24452 15976 24508
rect 15976 24452 15980 24508
rect 15916 24448 15980 24452
rect 45124 24508 45188 24512
rect 45124 24452 45128 24508
rect 45128 24452 45184 24508
rect 45184 24452 45188 24508
rect 45124 24448 45188 24452
rect 45204 24508 45268 24512
rect 45204 24452 45208 24508
rect 45208 24452 45264 24508
rect 45264 24452 45268 24508
rect 45204 24448 45268 24452
rect 45284 24508 45348 24512
rect 45284 24452 45288 24508
rect 45288 24452 45344 24508
rect 45344 24452 45348 24508
rect 45284 24448 45348 24452
rect 45364 24508 45428 24512
rect 45364 24452 45368 24508
rect 45368 24452 45424 24508
rect 45424 24452 45428 24508
rect 45364 24448 45428 24452
rect 74572 24508 74636 24512
rect 74572 24452 74576 24508
rect 74576 24452 74632 24508
rect 74632 24452 74636 24508
rect 74572 24448 74636 24452
rect 74652 24508 74716 24512
rect 74652 24452 74656 24508
rect 74656 24452 74712 24508
rect 74712 24452 74716 24508
rect 74652 24448 74716 24452
rect 74732 24508 74796 24512
rect 74732 24452 74736 24508
rect 74736 24452 74792 24508
rect 74792 24452 74796 24508
rect 74732 24448 74796 24452
rect 74812 24508 74876 24512
rect 74812 24452 74816 24508
rect 74816 24452 74872 24508
rect 74872 24452 74876 24508
rect 74812 24448 74876 24452
rect 104020 24508 104084 24512
rect 104020 24452 104024 24508
rect 104024 24452 104080 24508
rect 104080 24452 104084 24508
rect 104020 24448 104084 24452
rect 104100 24508 104164 24512
rect 104100 24452 104104 24508
rect 104104 24452 104160 24508
rect 104160 24452 104164 24508
rect 104100 24448 104164 24452
rect 104180 24508 104244 24512
rect 104180 24452 104184 24508
rect 104184 24452 104240 24508
rect 104240 24452 104244 24508
rect 104180 24448 104244 24452
rect 104260 24508 104324 24512
rect 104260 24452 104264 24508
rect 104264 24452 104320 24508
rect 104320 24452 104324 24508
rect 104260 24448 104324 24452
rect 30400 23964 30464 23968
rect 30400 23908 30404 23964
rect 30404 23908 30460 23964
rect 30460 23908 30464 23964
rect 30400 23904 30464 23908
rect 30480 23964 30544 23968
rect 30480 23908 30484 23964
rect 30484 23908 30540 23964
rect 30540 23908 30544 23964
rect 30480 23904 30544 23908
rect 30560 23964 30624 23968
rect 30560 23908 30564 23964
rect 30564 23908 30620 23964
rect 30620 23908 30624 23964
rect 30560 23904 30624 23908
rect 30640 23964 30704 23968
rect 30640 23908 30644 23964
rect 30644 23908 30700 23964
rect 30700 23908 30704 23964
rect 30640 23904 30704 23908
rect 59848 23964 59912 23968
rect 59848 23908 59852 23964
rect 59852 23908 59908 23964
rect 59908 23908 59912 23964
rect 59848 23904 59912 23908
rect 59928 23964 59992 23968
rect 59928 23908 59932 23964
rect 59932 23908 59988 23964
rect 59988 23908 59992 23964
rect 59928 23904 59992 23908
rect 60008 23964 60072 23968
rect 60008 23908 60012 23964
rect 60012 23908 60068 23964
rect 60068 23908 60072 23964
rect 60008 23904 60072 23908
rect 60088 23964 60152 23968
rect 60088 23908 60092 23964
rect 60092 23908 60148 23964
rect 60148 23908 60152 23964
rect 60088 23904 60152 23908
rect 89296 23964 89360 23968
rect 89296 23908 89300 23964
rect 89300 23908 89356 23964
rect 89356 23908 89360 23964
rect 89296 23904 89360 23908
rect 89376 23964 89440 23968
rect 89376 23908 89380 23964
rect 89380 23908 89436 23964
rect 89436 23908 89440 23964
rect 89376 23904 89440 23908
rect 89456 23964 89520 23968
rect 89456 23908 89460 23964
rect 89460 23908 89516 23964
rect 89516 23908 89520 23964
rect 89456 23904 89520 23908
rect 89536 23964 89600 23968
rect 89536 23908 89540 23964
rect 89540 23908 89596 23964
rect 89596 23908 89600 23964
rect 89536 23904 89600 23908
rect 15676 23420 15740 23424
rect 15676 23364 15680 23420
rect 15680 23364 15736 23420
rect 15736 23364 15740 23420
rect 15676 23360 15740 23364
rect 15756 23420 15820 23424
rect 15756 23364 15760 23420
rect 15760 23364 15816 23420
rect 15816 23364 15820 23420
rect 15756 23360 15820 23364
rect 15836 23420 15900 23424
rect 15836 23364 15840 23420
rect 15840 23364 15896 23420
rect 15896 23364 15900 23420
rect 15836 23360 15900 23364
rect 15916 23420 15980 23424
rect 15916 23364 15920 23420
rect 15920 23364 15976 23420
rect 15976 23364 15980 23420
rect 15916 23360 15980 23364
rect 45124 23420 45188 23424
rect 45124 23364 45128 23420
rect 45128 23364 45184 23420
rect 45184 23364 45188 23420
rect 45124 23360 45188 23364
rect 45204 23420 45268 23424
rect 45204 23364 45208 23420
rect 45208 23364 45264 23420
rect 45264 23364 45268 23420
rect 45204 23360 45268 23364
rect 45284 23420 45348 23424
rect 45284 23364 45288 23420
rect 45288 23364 45344 23420
rect 45344 23364 45348 23420
rect 45284 23360 45348 23364
rect 45364 23420 45428 23424
rect 45364 23364 45368 23420
rect 45368 23364 45424 23420
rect 45424 23364 45428 23420
rect 45364 23360 45428 23364
rect 74572 23420 74636 23424
rect 74572 23364 74576 23420
rect 74576 23364 74632 23420
rect 74632 23364 74636 23420
rect 74572 23360 74636 23364
rect 74652 23420 74716 23424
rect 74652 23364 74656 23420
rect 74656 23364 74712 23420
rect 74712 23364 74716 23420
rect 74652 23360 74716 23364
rect 74732 23420 74796 23424
rect 74732 23364 74736 23420
rect 74736 23364 74792 23420
rect 74792 23364 74796 23420
rect 74732 23360 74796 23364
rect 74812 23420 74876 23424
rect 74812 23364 74816 23420
rect 74816 23364 74872 23420
rect 74872 23364 74876 23420
rect 74812 23360 74876 23364
rect 104020 23420 104084 23424
rect 104020 23364 104024 23420
rect 104024 23364 104080 23420
rect 104080 23364 104084 23420
rect 104020 23360 104084 23364
rect 104100 23420 104164 23424
rect 104100 23364 104104 23420
rect 104104 23364 104160 23420
rect 104160 23364 104164 23420
rect 104100 23360 104164 23364
rect 104180 23420 104244 23424
rect 104180 23364 104184 23420
rect 104184 23364 104240 23420
rect 104240 23364 104244 23420
rect 104180 23360 104244 23364
rect 104260 23420 104324 23424
rect 104260 23364 104264 23420
rect 104264 23364 104320 23420
rect 104320 23364 104324 23420
rect 104260 23360 104324 23364
rect 30400 22876 30464 22880
rect 30400 22820 30404 22876
rect 30404 22820 30460 22876
rect 30460 22820 30464 22876
rect 30400 22816 30464 22820
rect 30480 22876 30544 22880
rect 30480 22820 30484 22876
rect 30484 22820 30540 22876
rect 30540 22820 30544 22876
rect 30480 22816 30544 22820
rect 30560 22876 30624 22880
rect 30560 22820 30564 22876
rect 30564 22820 30620 22876
rect 30620 22820 30624 22876
rect 30560 22816 30624 22820
rect 30640 22876 30704 22880
rect 30640 22820 30644 22876
rect 30644 22820 30700 22876
rect 30700 22820 30704 22876
rect 30640 22816 30704 22820
rect 59848 22876 59912 22880
rect 59848 22820 59852 22876
rect 59852 22820 59908 22876
rect 59908 22820 59912 22876
rect 59848 22816 59912 22820
rect 59928 22876 59992 22880
rect 59928 22820 59932 22876
rect 59932 22820 59988 22876
rect 59988 22820 59992 22876
rect 59928 22816 59992 22820
rect 60008 22876 60072 22880
rect 60008 22820 60012 22876
rect 60012 22820 60068 22876
rect 60068 22820 60072 22876
rect 60008 22816 60072 22820
rect 60088 22876 60152 22880
rect 60088 22820 60092 22876
rect 60092 22820 60148 22876
rect 60148 22820 60152 22876
rect 60088 22816 60152 22820
rect 89296 22876 89360 22880
rect 89296 22820 89300 22876
rect 89300 22820 89356 22876
rect 89356 22820 89360 22876
rect 89296 22816 89360 22820
rect 89376 22876 89440 22880
rect 89376 22820 89380 22876
rect 89380 22820 89436 22876
rect 89436 22820 89440 22876
rect 89376 22816 89440 22820
rect 89456 22876 89520 22880
rect 89456 22820 89460 22876
rect 89460 22820 89516 22876
rect 89516 22820 89520 22876
rect 89456 22816 89520 22820
rect 89536 22876 89600 22880
rect 89536 22820 89540 22876
rect 89540 22820 89596 22876
rect 89596 22820 89600 22876
rect 89536 22816 89600 22820
rect 15676 22332 15740 22336
rect 15676 22276 15680 22332
rect 15680 22276 15736 22332
rect 15736 22276 15740 22332
rect 15676 22272 15740 22276
rect 15756 22332 15820 22336
rect 15756 22276 15760 22332
rect 15760 22276 15816 22332
rect 15816 22276 15820 22332
rect 15756 22272 15820 22276
rect 15836 22332 15900 22336
rect 15836 22276 15840 22332
rect 15840 22276 15896 22332
rect 15896 22276 15900 22332
rect 15836 22272 15900 22276
rect 15916 22332 15980 22336
rect 15916 22276 15920 22332
rect 15920 22276 15976 22332
rect 15976 22276 15980 22332
rect 15916 22272 15980 22276
rect 45124 22332 45188 22336
rect 45124 22276 45128 22332
rect 45128 22276 45184 22332
rect 45184 22276 45188 22332
rect 45124 22272 45188 22276
rect 45204 22332 45268 22336
rect 45204 22276 45208 22332
rect 45208 22276 45264 22332
rect 45264 22276 45268 22332
rect 45204 22272 45268 22276
rect 45284 22332 45348 22336
rect 45284 22276 45288 22332
rect 45288 22276 45344 22332
rect 45344 22276 45348 22332
rect 45284 22272 45348 22276
rect 45364 22332 45428 22336
rect 45364 22276 45368 22332
rect 45368 22276 45424 22332
rect 45424 22276 45428 22332
rect 45364 22272 45428 22276
rect 74572 22332 74636 22336
rect 74572 22276 74576 22332
rect 74576 22276 74632 22332
rect 74632 22276 74636 22332
rect 74572 22272 74636 22276
rect 74652 22332 74716 22336
rect 74652 22276 74656 22332
rect 74656 22276 74712 22332
rect 74712 22276 74716 22332
rect 74652 22272 74716 22276
rect 74732 22332 74796 22336
rect 74732 22276 74736 22332
rect 74736 22276 74792 22332
rect 74792 22276 74796 22332
rect 74732 22272 74796 22276
rect 74812 22332 74876 22336
rect 74812 22276 74816 22332
rect 74816 22276 74872 22332
rect 74872 22276 74876 22332
rect 74812 22272 74876 22276
rect 104020 22332 104084 22336
rect 104020 22276 104024 22332
rect 104024 22276 104080 22332
rect 104080 22276 104084 22332
rect 104020 22272 104084 22276
rect 104100 22332 104164 22336
rect 104100 22276 104104 22332
rect 104104 22276 104160 22332
rect 104160 22276 104164 22332
rect 104100 22272 104164 22276
rect 104180 22332 104244 22336
rect 104180 22276 104184 22332
rect 104184 22276 104240 22332
rect 104240 22276 104244 22332
rect 104180 22272 104244 22276
rect 104260 22332 104324 22336
rect 104260 22276 104264 22332
rect 104264 22276 104320 22332
rect 104320 22276 104324 22332
rect 104260 22272 104324 22276
rect 30400 21788 30464 21792
rect 30400 21732 30404 21788
rect 30404 21732 30460 21788
rect 30460 21732 30464 21788
rect 30400 21728 30464 21732
rect 30480 21788 30544 21792
rect 30480 21732 30484 21788
rect 30484 21732 30540 21788
rect 30540 21732 30544 21788
rect 30480 21728 30544 21732
rect 30560 21788 30624 21792
rect 30560 21732 30564 21788
rect 30564 21732 30620 21788
rect 30620 21732 30624 21788
rect 30560 21728 30624 21732
rect 30640 21788 30704 21792
rect 30640 21732 30644 21788
rect 30644 21732 30700 21788
rect 30700 21732 30704 21788
rect 30640 21728 30704 21732
rect 59848 21788 59912 21792
rect 59848 21732 59852 21788
rect 59852 21732 59908 21788
rect 59908 21732 59912 21788
rect 59848 21728 59912 21732
rect 59928 21788 59992 21792
rect 59928 21732 59932 21788
rect 59932 21732 59988 21788
rect 59988 21732 59992 21788
rect 59928 21728 59992 21732
rect 60008 21788 60072 21792
rect 60008 21732 60012 21788
rect 60012 21732 60068 21788
rect 60068 21732 60072 21788
rect 60008 21728 60072 21732
rect 60088 21788 60152 21792
rect 60088 21732 60092 21788
rect 60092 21732 60148 21788
rect 60148 21732 60152 21788
rect 60088 21728 60152 21732
rect 89296 21788 89360 21792
rect 89296 21732 89300 21788
rect 89300 21732 89356 21788
rect 89356 21732 89360 21788
rect 89296 21728 89360 21732
rect 89376 21788 89440 21792
rect 89376 21732 89380 21788
rect 89380 21732 89436 21788
rect 89436 21732 89440 21788
rect 89376 21728 89440 21732
rect 89456 21788 89520 21792
rect 89456 21732 89460 21788
rect 89460 21732 89516 21788
rect 89516 21732 89520 21788
rect 89456 21728 89520 21732
rect 89536 21788 89600 21792
rect 89536 21732 89540 21788
rect 89540 21732 89596 21788
rect 89596 21732 89600 21788
rect 89536 21728 89600 21732
rect 15676 21244 15740 21248
rect 15676 21188 15680 21244
rect 15680 21188 15736 21244
rect 15736 21188 15740 21244
rect 15676 21184 15740 21188
rect 15756 21244 15820 21248
rect 15756 21188 15760 21244
rect 15760 21188 15816 21244
rect 15816 21188 15820 21244
rect 15756 21184 15820 21188
rect 15836 21244 15900 21248
rect 15836 21188 15840 21244
rect 15840 21188 15896 21244
rect 15896 21188 15900 21244
rect 15836 21184 15900 21188
rect 15916 21244 15980 21248
rect 15916 21188 15920 21244
rect 15920 21188 15976 21244
rect 15976 21188 15980 21244
rect 15916 21184 15980 21188
rect 45124 21244 45188 21248
rect 45124 21188 45128 21244
rect 45128 21188 45184 21244
rect 45184 21188 45188 21244
rect 45124 21184 45188 21188
rect 45204 21244 45268 21248
rect 45204 21188 45208 21244
rect 45208 21188 45264 21244
rect 45264 21188 45268 21244
rect 45204 21184 45268 21188
rect 45284 21244 45348 21248
rect 45284 21188 45288 21244
rect 45288 21188 45344 21244
rect 45344 21188 45348 21244
rect 45284 21184 45348 21188
rect 45364 21244 45428 21248
rect 45364 21188 45368 21244
rect 45368 21188 45424 21244
rect 45424 21188 45428 21244
rect 45364 21184 45428 21188
rect 74572 21244 74636 21248
rect 74572 21188 74576 21244
rect 74576 21188 74632 21244
rect 74632 21188 74636 21244
rect 74572 21184 74636 21188
rect 74652 21244 74716 21248
rect 74652 21188 74656 21244
rect 74656 21188 74712 21244
rect 74712 21188 74716 21244
rect 74652 21184 74716 21188
rect 74732 21244 74796 21248
rect 74732 21188 74736 21244
rect 74736 21188 74792 21244
rect 74792 21188 74796 21244
rect 74732 21184 74796 21188
rect 74812 21244 74876 21248
rect 74812 21188 74816 21244
rect 74816 21188 74872 21244
rect 74872 21188 74876 21244
rect 74812 21184 74876 21188
rect 104020 21244 104084 21248
rect 104020 21188 104024 21244
rect 104024 21188 104080 21244
rect 104080 21188 104084 21244
rect 104020 21184 104084 21188
rect 104100 21244 104164 21248
rect 104100 21188 104104 21244
rect 104104 21188 104160 21244
rect 104160 21188 104164 21244
rect 104100 21184 104164 21188
rect 104180 21244 104244 21248
rect 104180 21188 104184 21244
rect 104184 21188 104240 21244
rect 104240 21188 104244 21244
rect 104180 21184 104244 21188
rect 104260 21244 104324 21248
rect 104260 21188 104264 21244
rect 104264 21188 104320 21244
rect 104320 21188 104324 21244
rect 104260 21184 104324 21188
rect 30400 20700 30464 20704
rect 30400 20644 30404 20700
rect 30404 20644 30460 20700
rect 30460 20644 30464 20700
rect 30400 20640 30464 20644
rect 30480 20700 30544 20704
rect 30480 20644 30484 20700
rect 30484 20644 30540 20700
rect 30540 20644 30544 20700
rect 30480 20640 30544 20644
rect 30560 20700 30624 20704
rect 30560 20644 30564 20700
rect 30564 20644 30620 20700
rect 30620 20644 30624 20700
rect 30560 20640 30624 20644
rect 30640 20700 30704 20704
rect 30640 20644 30644 20700
rect 30644 20644 30700 20700
rect 30700 20644 30704 20700
rect 30640 20640 30704 20644
rect 59848 20700 59912 20704
rect 59848 20644 59852 20700
rect 59852 20644 59908 20700
rect 59908 20644 59912 20700
rect 59848 20640 59912 20644
rect 59928 20700 59992 20704
rect 59928 20644 59932 20700
rect 59932 20644 59988 20700
rect 59988 20644 59992 20700
rect 59928 20640 59992 20644
rect 60008 20700 60072 20704
rect 60008 20644 60012 20700
rect 60012 20644 60068 20700
rect 60068 20644 60072 20700
rect 60008 20640 60072 20644
rect 60088 20700 60152 20704
rect 60088 20644 60092 20700
rect 60092 20644 60148 20700
rect 60148 20644 60152 20700
rect 60088 20640 60152 20644
rect 89296 20700 89360 20704
rect 89296 20644 89300 20700
rect 89300 20644 89356 20700
rect 89356 20644 89360 20700
rect 89296 20640 89360 20644
rect 89376 20700 89440 20704
rect 89376 20644 89380 20700
rect 89380 20644 89436 20700
rect 89436 20644 89440 20700
rect 89376 20640 89440 20644
rect 89456 20700 89520 20704
rect 89456 20644 89460 20700
rect 89460 20644 89516 20700
rect 89516 20644 89520 20700
rect 89456 20640 89520 20644
rect 89536 20700 89600 20704
rect 89536 20644 89540 20700
rect 89540 20644 89596 20700
rect 89596 20644 89600 20700
rect 89536 20640 89600 20644
rect 15676 20156 15740 20160
rect 15676 20100 15680 20156
rect 15680 20100 15736 20156
rect 15736 20100 15740 20156
rect 15676 20096 15740 20100
rect 15756 20156 15820 20160
rect 15756 20100 15760 20156
rect 15760 20100 15816 20156
rect 15816 20100 15820 20156
rect 15756 20096 15820 20100
rect 15836 20156 15900 20160
rect 15836 20100 15840 20156
rect 15840 20100 15896 20156
rect 15896 20100 15900 20156
rect 15836 20096 15900 20100
rect 15916 20156 15980 20160
rect 15916 20100 15920 20156
rect 15920 20100 15976 20156
rect 15976 20100 15980 20156
rect 15916 20096 15980 20100
rect 45124 20156 45188 20160
rect 45124 20100 45128 20156
rect 45128 20100 45184 20156
rect 45184 20100 45188 20156
rect 45124 20096 45188 20100
rect 45204 20156 45268 20160
rect 45204 20100 45208 20156
rect 45208 20100 45264 20156
rect 45264 20100 45268 20156
rect 45204 20096 45268 20100
rect 45284 20156 45348 20160
rect 45284 20100 45288 20156
rect 45288 20100 45344 20156
rect 45344 20100 45348 20156
rect 45284 20096 45348 20100
rect 45364 20156 45428 20160
rect 45364 20100 45368 20156
rect 45368 20100 45424 20156
rect 45424 20100 45428 20156
rect 45364 20096 45428 20100
rect 74572 20156 74636 20160
rect 74572 20100 74576 20156
rect 74576 20100 74632 20156
rect 74632 20100 74636 20156
rect 74572 20096 74636 20100
rect 74652 20156 74716 20160
rect 74652 20100 74656 20156
rect 74656 20100 74712 20156
rect 74712 20100 74716 20156
rect 74652 20096 74716 20100
rect 74732 20156 74796 20160
rect 74732 20100 74736 20156
rect 74736 20100 74792 20156
rect 74792 20100 74796 20156
rect 74732 20096 74796 20100
rect 74812 20156 74876 20160
rect 74812 20100 74816 20156
rect 74816 20100 74872 20156
rect 74872 20100 74876 20156
rect 74812 20096 74876 20100
rect 104020 20156 104084 20160
rect 104020 20100 104024 20156
rect 104024 20100 104080 20156
rect 104080 20100 104084 20156
rect 104020 20096 104084 20100
rect 104100 20156 104164 20160
rect 104100 20100 104104 20156
rect 104104 20100 104160 20156
rect 104160 20100 104164 20156
rect 104100 20096 104164 20100
rect 104180 20156 104244 20160
rect 104180 20100 104184 20156
rect 104184 20100 104240 20156
rect 104240 20100 104244 20156
rect 104180 20096 104244 20100
rect 104260 20156 104324 20160
rect 104260 20100 104264 20156
rect 104264 20100 104320 20156
rect 104320 20100 104324 20156
rect 104260 20096 104324 20100
rect 30400 19612 30464 19616
rect 30400 19556 30404 19612
rect 30404 19556 30460 19612
rect 30460 19556 30464 19612
rect 30400 19552 30464 19556
rect 30480 19612 30544 19616
rect 30480 19556 30484 19612
rect 30484 19556 30540 19612
rect 30540 19556 30544 19612
rect 30480 19552 30544 19556
rect 30560 19612 30624 19616
rect 30560 19556 30564 19612
rect 30564 19556 30620 19612
rect 30620 19556 30624 19612
rect 30560 19552 30624 19556
rect 30640 19612 30704 19616
rect 30640 19556 30644 19612
rect 30644 19556 30700 19612
rect 30700 19556 30704 19612
rect 30640 19552 30704 19556
rect 59848 19612 59912 19616
rect 59848 19556 59852 19612
rect 59852 19556 59908 19612
rect 59908 19556 59912 19612
rect 59848 19552 59912 19556
rect 59928 19612 59992 19616
rect 59928 19556 59932 19612
rect 59932 19556 59988 19612
rect 59988 19556 59992 19612
rect 59928 19552 59992 19556
rect 60008 19612 60072 19616
rect 60008 19556 60012 19612
rect 60012 19556 60068 19612
rect 60068 19556 60072 19612
rect 60008 19552 60072 19556
rect 60088 19612 60152 19616
rect 60088 19556 60092 19612
rect 60092 19556 60148 19612
rect 60148 19556 60152 19612
rect 60088 19552 60152 19556
rect 89296 19612 89360 19616
rect 89296 19556 89300 19612
rect 89300 19556 89356 19612
rect 89356 19556 89360 19612
rect 89296 19552 89360 19556
rect 89376 19612 89440 19616
rect 89376 19556 89380 19612
rect 89380 19556 89436 19612
rect 89436 19556 89440 19612
rect 89376 19552 89440 19556
rect 89456 19612 89520 19616
rect 89456 19556 89460 19612
rect 89460 19556 89516 19612
rect 89516 19556 89520 19612
rect 89456 19552 89520 19556
rect 89536 19612 89600 19616
rect 89536 19556 89540 19612
rect 89540 19556 89596 19612
rect 89596 19556 89600 19612
rect 89536 19552 89600 19556
rect 15676 19068 15740 19072
rect 15676 19012 15680 19068
rect 15680 19012 15736 19068
rect 15736 19012 15740 19068
rect 15676 19008 15740 19012
rect 15756 19068 15820 19072
rect 15756 19012 15760 19068
rect 15760 19012 15816 19068
rect 15816 19012 15820 19068
rect 15756 19008 15820 19012
rect 15836 19068 15900 19072
rect 15836 19012 15840 19068
rect 15840 19012 15896 19068
rect 15896 19012 15900 19068
rect 15836 19008 15900 19012
rect 15916 19068 15980 19072
rect 15916 19012 15920 19068
rect 15920 19012 15976 19068
rect 15976 19012 15980 19068
rect 15916 19008 15980 19012
rect 45124 19068 45188 19072
rect 45124 19012 45128 19068
rect 45128 19012 45184 19068
rect 45184 19012 45188 19068
rect 45124 19008 45188 19012
rect 45204 19068 45268 19072
rect 45204 19012 45208 19068
rect 45208 19012 45264 19068
rect 45264 19012 45268 19068
rect 45204 19008 45268 19012
rect 45284 19068 45348 19072
rect 45284 19012 45288 19068
rect 45288 19012 45344 19068
rect 45344 19012 45348 19068
rect 45284 19008 45348 19012
rect 45364 19068 45428 19072
rect 45364 19012 45368 19068
rect 45368 19012 45424 19068
rect 45424 19012 45428 19068
rect 45364 19008 45428 19012
rect 74572 19068 74636 19072
rect 74572 19012 74576 19068
rect 74576 19012 74632 19068
rect 74632 19012 74636 19068
rect 74572 19008 74636 19012
rect 74652 19068 74716 19072
rect 74652 19012 74656 19068
rect 74656 19012 74712 19068
rect 74712 19012 74716 19068
rect 74652 19008 74716 19012
rect 74732 19068 74796 19072
rect 74732 19012 74736 19068
rect 74736 19012 74792 19068
rect 74792 19012 74796 19068
rect 74732 19008 74796 19012
rect 74812 19068 74876 19072
rect 74812 19012 74816 19068
rect 74816 19012 74872 19068
rect 74872 19012 74876 19068
rect 74812 19008 74876 19012
rect 104020 19068 104084 19072
rect 104020 19012 104024 19068
rect 104024 19012 104080 19068
rect 104080 19012 104084 19068
rect 104020 19008 104084 19012
rect 104100 19068 104164 19072
rect 104100 19012 104104 19068
rect 104104 19012 104160 19068
rect 104160 19012 104164 19068
rect 104100 19008 104164 19012
rect 104180 19068 104244 19072
rect 104180 19012 104184 19068
rect 104184 19012 104240 19068
rect 104240 19012 104244 19068
rect 104180 19008 104244 19012
rect 104260 19068 104324 19072
rect 104260 19012 104264 19068
rect 104264 19012 104320 19068
rect 104320 19012 104324 19068
rect 104260 19008 104324 19012
rect 30400 18524 30464 18528
rect 30400 18468 30404 18524
rect 30404 18468 30460 18524
rect 30460 18468 30464 18524
rect 30400 18464 30464 18468
rect 30480 18524 30544 18528
rect 30480 18468 30484 18524
rect 30484 18468 30540 18524
rect 30540 18468 30544 18524
rect 30480 18464 30544 18468
rect 30560 18524 30624 18528
rect 30560 18468 30564 18524
rect 30564 18468 30620 18524
rect 30620 18468 30624 18524
rect 30560 18464 30624 18468
rect 30640 18524 30704 18528
rect 30640 18468 30644 18524
rect 30644 18468 30700 18524
rect 30700 18468 30704 18524
rect 30640 18464 30704 18468
rect 59848 18524 59912 18528
rect 59848 18468 59852 18524
rect 59852 18468 59908 18524
rect 59908 18468 59912 18524
rect 59848 18464 59912 18468
rect 59928 18524 59992 18528
rect 59928 18468 59932 18524
rect 59932 18468 59988 18524
rect 59988 18468 59992 18524
rect 59928 18464 59992 18468
rect 60008 18524 60072 18528
rect 60008 18468 60012 18524
rect 60012 18468 60068 18524
rect 60068 18468 60072 18524
rect 60008 18464 60072 18468
rect 60088 18524 60152 18528
rect 60088 18468 60092 18524
rect 60092 18468 60148 18524
rect 60148 18468 60152 18524
rect 60088 18464 60152 18468
rect 89296 18524 89360 18528
rect 89296 18468 89300 18524
rect 89300 18468 89356 18524
rect 89356 18468 89360 18524
rect 89296 18464 89360 18468
rect 89376 18524 89440 18528
rect 89376 18468 89380 18524
rect 89380 18468 89436 18524
rect 89436 18468 89440 18524
rect 89376 18464 89440 18468
rect 89456 18524 89520 18528
rect 89456 18468 89460 18524
rect 89460 18468 89516 18524
rect 89516 18468 89520 18524
rect 89456 18464 89520 18468
rect 89536 18524 89600 18528
rect 89536 18468 89540 18524
rect 89540 18468 89596 18524
rect 89596 18468 89600 18524
rect 89536 18464 89600 18468
rect 15676 17980 15740 17984
rect 15676 17924 15680 17980
rect 15680 17924 15736 17980
rect 15736 17924 15740 17980
rect 15676 17920 15740 17924
rect 15756 17980 15820 17984
rect 15756 17924 15760 17980
rect 15760 17924 15816 17980
rect 15816 17924 15820 17980
rect 15756 17920 15820 17924
rect 15836 17980 15900 17984
rect 15836 17924 15840 17980
rect 15840 17924 15896 17980
rect 15896 17924 15900 17980
rect 15836 17920 15900 17924
rect 15916 17980 15980 17984
rect 15916 17924 15920 17980
rect 15920 17924 15976 17980
rect 15976 17924 15980 17980
rect 15916 17920 15980 17924
rect 45124 17980 45188 17984
rect 45124 17924 45128 17980
rect 45128 17924 45184 17980
rect 45184 17924 45188 17980
rect 45124 17920 45188 17924
rect 45204 17980 45268 17984
rect 45204 17924 45208 17980
rect 45208 17924 45264 17980
rect 45264 17924 45268 17980
rect 45204 17920 45268 17924
rect 45284 17980 45348 17984
rect 45284 17924 45288 17980
rect 45288 17924 45344 17980
rect 45344 17924 45348 17980
rect 45284 17920 45348 17924
rect 45364 17980 45428 17984
rect 45364 17924 45368 17980
rect 45368 17924 45424 17980
rect 45424 17924 45428 17980
rect 45364 17920 45428 17924
rect 74572 17980 74636 17984
rect 74572 17924 74576 17980
rect 74576 17924 74632 17980
rect 74632 17924 74636 17980
rect 74572 17920 74636 17924
rect 74652 17980 74716 17984
rect 74652 17924 74656 17980
rect 74656 17924 74712 17980
rect 74712 17924 74716 17980
rect 74652 17920 74716 17924
rect 74732 17980 74796 17984
rect 74732 17924 74736 17980
rect 74736 17924 74792 17980
rect 74792 17924 74796 17980
rect 74732 17920 74796 17924
rect 74812 17980 74876 17984
rect 74812 17924 74816 17980
rect 74816 17924 74872 17980
rect 74872 17924 74876 17980
rect 74812 17920 74876 17924
rect 104020 17980 104084 17984
rect 104020 17924 104024 17980
rect 104024 17924 104080 17980
rect 104080 17924 104084 17980
rect 104020 17920 104084 17924
rect 104100 17980 104164 17984
rect 104100 17924 104104 17980
rect 104104 17924 104160 17980
rect 104160 17924 104164 17980
rect 104100 17920 104164 17924
rect 104180 17980 104244 17984
rect 104180 17924 104184 17980
rect 104184 17924 104240 17980
rect 104240 17924 104244 17980
rect 104180 17920 104244 17924
rect 104260 17980 104324 17984
rect 104260 17924 104264 17980
rect 104264 17924 104320 17980
rect 104320 17924 104324 17980
rect 104260 17920 104324 17924
rect 30400 17436 30464 17440
rect 30400 17380 30404 17436
rect 30404 17380 30460 17436
rect 30460 17380 30464 17436
rect 30400 17376 30464 17380
rect 30480 17436 30544 17440
rect 30480 17380 30484 17436
rect 30484 17380 30540 17436
rect 30540 17380 30544 17436
rect 30480 17376 30544 17380
rect 30560 17436 30624 17440
rect 30560 17380 30564 17436
rect 30564 17380 30620 17436
rect 30620 17380 30624 17436
rect 30560 17376 30624 17380
rect 30640 17436 30704 17440
rect 30640 17380 30644 17436
rect 30644 17380 30700 17436
rect 30700 17380 30704 17436
rect 30640 17376 30704 17380
rect 59848 17436 59912 17440
rect 59848 17380 59852 17436
rect 59852 17380 59908 17436
rect 59908 17380 59912 17436
rect 59848 17376 59912 17380
rect 59928 17436 59992 17440
rect 59928 17380 59932 17436
rect 59932 17380 59988 17436
rect 59988 17380 59992 17436
rect 59928 17376 59992 17380
rect 60008 17436 60072 17440
rect 60008 17380 60012 17436
rect 60012 17380 60068 17436
rect 60068 17380 60072 17436
rect 60008 17376 60072 17380
rect 60088 17436 60152 17440
rect 60088 17380 60092 17436
rect 60092 17380 60148 17436
rect 60148 17380 60152 17436
rect 60088 17376 60152 17380
rect 89296 17436 89360 17440
rect 89296 17380 89300 17436
rect 89300 17380 89356 17436
rect 89356 17380 89360 17436
rect 89296 17376 89360 17380
rect 89376 17436 89440 17440
rect 89376 17380 89380 17436
rect 89380 17380 89436 17436
rect 89436 17380 89440 17436
rect 89376 17376 89440 17380
rect 89456 17436 89520 17440
rect 89456 17380 89460 17436
rect 89460 17380 89516 17436
rect 89516 17380 89520 17436
rect 89456 17376 89520 17380
rect 89536 17436 89600 17440
rect 89536 17380 89540 17436
rect 89540 17380 89596 17436
rect 89596 17380 89600 17436
rect 89536 17376 89600 17380
rect 15676 16892 15740 16896
rect 15676 16836 15680 16892
rect 15680 16836 15736 16892
rect 15736 16836 15740 16892
rect 15676 16832 15740 16836
rect 15756 16892 15820 16896
rect 15756 16836 15760 16892
rect 15760 16836 15816 16892
rect 15816 16836 15820 16892
rect 15756 16832 15820 16836
rect 15836 16892 15900 16896
rect 15836 16836 15840 16892
rect 15840 16836 15896 16892
rect 15896 16836 15900 16892
rect 15836 16832 15900 16836
rect 15916 16892 15980 16896
rect 15916 16836 15920 16892
rect 15920 16836 15976 16892
rect 15976 16836 15980 16892
rect 15916 16832 15980 16836
rect 45124 16892 45188 16896
rect 45124 16836 45128 16892
rect 45128 16836 45184 16892
rect 45184 16836 45188 16892
rect 45124 16832 45188 16836
rect 45204 16892 45268 16896
rect 45204 16836 45208 16892
rect 45208 16836 45264 16892
rect 45264 16836 45268 16892
rect 45204 16832 45268 16836
rect 45284 16892 45348 16896
rect 45284 16836 45288 16892
rect 45288 16836 45344 16892
rect 45344 16836 45348 16892
rect 45284 16832 45348 16836
rect 45364 16892 45428 16896
rect 45364 16836 45368 16892
rect 45368 16836 45424 16892
rect 45424 16836 45428 16892
rect 45364 16832 45428 16836
rect 74572 16892 74636 16896
rect 74572 16836 74576 16892
rect 74576 16836 74632 16892
rect 74632 16836 74636 16892
rect 74572 16832 74636 16836
rect 74652 16892 74716 16896
rect 74652 16836 74656 16892
rect 74656 16836 74712 16892
rect 74712 16836 74716 16892
rect 74652 16832 74716 16836
rect 74732 16892 74796 16896
rect 74732 16836 74736 16892
rect 74736 16836 74792 16892
rect 74792 16836 74796 16892
rect 74732 16832 74796 16836
rect 74812 16892 74876 16896
rect 74812 16836 74816 16892
rect 74816 16836 74872 16892
rect 74872 16836 74876 16892
rect 74812 16832 74876 16836
rect 104020 16892 104084 16896
rect 104020 16836 104024 16892
rect 104024 16836 104080 16892
rect 104080 16836 104084 16892
rect 104020 16832 104084 16836
rect 104100 16892 104164 16896
rect 104100 16836 104104 16892
rect 104104 16836 104160 16892
rect 104160 16836 104164 16892
rect 104100 16832 104164 16836
rect 104180 16892 104244 16896
rect 104180 16836 104184 16892
rect 104184 16836 104240 16892
rect 104240 16836 104244 16892
rect 104180 16832 104244 16836
rect 104260 16892 104324 16896
rect 104260 16836 104264 16892
rect 104264 16836 104320 16892
rect 104320 16836 104324 16892
rect 104260 16832 104324 16836
rect 30400 16348 30464 16352
rect 30400 16292 30404 16348
rect 30404 16292 30460 16348
rect 30460 16292 30464 16348
rect 30400 16288 30464 16292
rect 30480 16348 30544 16352
rect 30480 16292 30484 16348
rect 30484 16292 30540 16348
rect 30540 16292 30544 16348
rect 30480 16288 30544 16292
rect 30560 16348 30624 16352
rect 30560 16292 30564 16348
rect 30564 16292 30620 16348
rect 30620 16292 30624 16348
rect 30560 16288 30624 16292
rect 30640 16348 30704 16352
rect 30640 16292 30644 16348
rect 30644 16292 30700 16348
rect 30700 16292 30704 16348
rect 30640 16288 30704 16292
rect 59848 16348 59912 16352
rect 59848 16292 59852 16348
rect 59852 16292 59908 16348
rect 59908 16292 59912 16348
rect 59848 16288 59912 16292
rect 59928 16348 59992 16352
rect 59928 16292 59932 16348
rect 59932 16292 59988 16348
rect 59988 16292 59992 16348
rect 59928 16288 59992 16292
rect 60008 16348 60072 16352
rect 60008 16292 60012 16348
rect 60012 16292 60068 16348
rect 60068 16292 60072 16348
rect 60008 16288 60072 16292
rect 60088 16348 60152 16352
rect 60088 16292 60092 16348
rect 60092 16292 60148 16348
rect 60148 16292 60152 16348
rect 60088 16288 60152 16292
rect 89296 16348 89360 16352
rect 89296 16292 89300 16348
rect 89300 16292 89356 16348
rect 89356 16292 89360 16348
rect 89296 16288 89360 16292
rect 89376 16348 89440 16352
rect 89376 16292 89380 16348
rect 89380 16292 89436 16348
rect 89436 16292 89440 16348
rect 89376 16288 89440 16292
rect 89456 16348 89520 16352
rect 89456 16292 89460 16348
rect 89460 16292 89516 16348
rect 89516 16292 89520 16348
rect 89456 16288 89520 16292
rect 89536 16348 89600 16352
rect 89536 16292 89540 16348
rect 89540 16292 89596 16348
rect 89596 16292 89600 16348
rect 89536 16288 89600 16292
rect 15676 15804 15740 15808
rect 15676 15748 15680 15804
rect 15680 15748 15736 15804
rect 15736 15748 15740 15804
rect 15676 15744 15740 15748
rect 15756 15804 15820 15808
rect 15756 15748 15760 15804
rect 15760 15748 15816 15804
rect 15816 15748 15820 15804
rect 15756 15744 15820 15748
rect 15836 15804 15900 15808
rect 15836 15748 15840 15804
rect 15840 15748 15896 15804
rect 15896 15748 15900 15804
rect 15836 15744 15900 15748
rect 15916 15804 15980 15808
rect 15916 15748 15920 15804
rect 15920 15748 15976 15804
rect 15976 15748 15980 15804
rect 15916 15744 15980 15748
rect 45124 15804 45188 15808
rect 45124 15748 45128 15804
rect 45128 15748 45184 15804
rect 45184 15748 45188 15804
rect 45124 15744 45188 15748
rect 45204 15804 45268 15808
rect 45204 15748 45208 15804
rect 45208 15748 45264 15804
rect 45264 15748 45268 15804
rect 45204 15744 45268 15748
rect 45284 15804 45348 15808
rect 45284 15748 45288 15804
rect 45288 15748 45344 15804
rect 45344 15748 45348 15804
rect 45284 15744 45348 15748
rect 45364 15804 45428 15808
rect 45364 15748 45368 15804
rect 45368 15748 45424 15804
rect 45424 15748 45428 15804
rect 45364 15744 45428 15748
rect 74572 15804 74636 15808
rect 74572 15748 74576 15804
rect 74576 15748 74632 15804
rect 74632 15748 74636 15804
rect 74572 15744 74636 15748
rect 74652 15804 74716 15808
rect 74652 15748 74656 15804
rect 74656 15748 74712 15804
rect 74712 15748 74716 15804
rect 74652 15744 74716 15748
rect 74732 15804 74796 15808
rect 74732 15748 74736 15804
rect 74736 15748 74792 15804
rect 74792 15748 74796 15804
rect 74732 15744 74796 15748
rect 74812 15804 74876 15808
rect 74812 15748 74816 15804
rect 74816 15748 74872 15804
rect 74872 15748 74876 15804
rect 74812 15744 74876 15748
rect 104020 15804 104084 15808
rect 104020 15748 104024 15804
rect 104024 15748 104080 15804
rect 104080 15748 104084 15804
rect 104020 15744 104084 15748
rect 104100 15804 104164 15808
rect 104100 15748 104104 15804
rect 104104 15748 104160 15804
rect 104160 15748 104164 15804
rect 104100 15744 104164 15748
rect 104180 15804 104244 15808
rect 104180 15748 104184 15804
rect 104184 15748 104240 15804
rect 104240 15748 104244 15804
rect 104180 15744 104244 15748
rect 104260 15804 104324 15808
rect 104260 15748 104264 15804
rect 104264 15748 104320 15804
rect 104320 15748 104324 15804
rect 104260 15744 104324 15748
rect 30400 15260 30464 15264
rect 30400 15204 30404 15260
rect 30404 15204 30460 15260
rect 30460 15204 30464 15260
rect 30400 15200 30464 15204
rect 30480 15260 30544 15264
rect 30480 15204 30484 15260
rect 30484 15204 30540 15260
rect 30540 15204 30544 15260
rect 30480 15200 30544 15204
rect 30560 15260 30624 15264
rect 30560 15204 30564 15260
rect 30564 15204 30620 15260
rect 30620 15204 30624 15260
rect 30560 15200 30624 15204
rect 30640 15260 30704 15264
rect 30640 15204 30644 15260
rect 30644 15204 30700 15260
rect 30700 15204 30704 15260
rect 30640 15200 30704 15204
rect 59848 15260 59912 15264
rect 59848 15204 59852 15260
rect 59852 15204 59908 15260
rect 59908 15204 59912 15260
rect 59848 15200 59912 15204
rect 59928 15260 59992 15264
rect 59928 15204 59932 15260
rect 59932 15204 59988 15260
rect 59988 15204 59992 15260
rect 59928 15200 59992 15204
rect 60008 15260 60072 15264
rect 60008 15204 60012 15260
rect 60012 15204 60068 15260
rect 60068 15204 60072 15260
rect 60008 15200 60072 15204
rect 60088 15260 60152 15264
rect 60088 15204 60092 15260
rect 60092 15204 60148 15260
rect 60148 15204 60152 15260
rect 60088 15200 60152 15204
rect 89296 15260 89360 15264
rect 89296 15204 89300 15260
rect 89300 15204 89356 15260
rect 89356 15204 89360 15260
rect 89296 15200 89360 15204
rect 89376 15260 89440 15264
rect 89376 15204 89380 15260
rect 89380 15204 89436 15260
rect 89436 15204 89440 15260
rect 89376 15200 89440 15204
rect 89456 15260 89520 15264
rect 89456 15204 89460 15260
rect 89460 15204 89516 15260
rect 89516 15204 89520 15260
rect 89456 15200 89520 15204
rect 89536 15260 89600 15264
rect 89536 15204 89540 15260
rect 89540 15204 89596 15260
rect 89596 15204 89600 15260
rect 89536 15200 89600 15204
rect 15676 14716 15740 14720
rect 15676 14660 15680 14716
rect 15680 14660 15736 14716
rect 15736 14660 15740 14716
rect 15676 14656 15740 14660
rect 15756 14716 15820 14720
rect 15756 14660 15760 14716
rect 15760 14660 15816 14716
rect 15816 14660 15820 14716
rect 15756 14656 15820 14660
rect 15836 14716 15900 14720
rect 15836 14660 15840 14716
rect 15840 14660 15896 14716
rect 15896 14660 15900 14716
rect 15836 14656 15900 14660
rect 15916 14716 15980 14720
rect 15916 14660 15920 14716
rect 15920 14660 15976 14716
rect 15976 14660 15980 14716
rect 15916 14656 15980 14660
rect 45124 14716 45188 14720
rect 45124 14660 45128 14716
rect 45128 14660 45184 14716
rect 45184 14660 45188 14716
rect 45124 14656 45188 14660
rect 45204 14716 45268 14720
rect 45204 14660 45208 14716
rect 45208 14660 45264 14716
rect 45264 14660 45268 14716
rect 45204 14656 45268 14660
rect 45284 14716 45348 14720
rect 45284 14660 45288 14716
rect 45288 14660 45344 14716
rect 45344 14660 45348 14716
rect 45284 14656 45348 14660
rect 45364 14716 45428 14720
rect 45364 14660 45368 14716
rect 45368 14660 45424 14716
rect 45424 14660 45428 14716
rect 45364 14656 45428 14660
rect 74572 14716 74636 14720
rect 74572 14660 74576 14716
rect 74576 14660 74632 14716
rect 74632 14660 74636 14716
rect 74572 14656 74636 14660
rect 74652 14716 74716 14720
rect 74652 14660 74656 14716
rect 74656 14660 74712 14716
rect 74712 14660 74716 14716
rect 74652 14656 74716 14660
rect 74732 14716 74796 14720
rect 74732 14660 74736 14716
rect 74736 14660 74792 14716
rect 74792 14660 74796 14716
rect 74732 14656 74796 14660
rect 74812 14716 74876 14720
rect 74812 14660 74816 14716
rect 74816 14660 74872 14716
rect 74872 14660 74876 14716
rect 74812 14656 74876 14660
rect 104020 14716 104084 14720
rect 104020 14660 104024 14716
rect 104024 14660 104080 14716
rect 104080 14660 104084 14716
rect 104020 14656 104084 14660
rect 104100 14716 104164 14720
rect 104100 14660 104104 14716
rect 104104 14660 104160 14716
rect 104160 14660 104164 14716
rect 104100 14656 104164 14660
rect 104180 14716 104244 14720
rect 104180 14660 104184 14716
rect 104184 14660 104240 14716
rect 104240 14660 104244 14716
rect 104180 14656 104244 14660
rect 104260 14716 104324 14720
rect 104260 14660 104264 14716
rect 104264 14660 104320 14716
rect 104320 14660 104324 14716
rect 104260 14656 104324 14660
rect 30400 14172 30464 14176
rect 30400 14116 30404 14172
rect 30404 14116 30460 14172
rect 30460 14116 30464 14172
rect 30400 14112 30464 14116
rect 30480 14172 30544 14176
rect 30480 14116 30484 14172
rect 30484 14116 30540 14172
rect 30540 14116 30544 14172
rect 30480 14112 30544 14116
rect 30560 14172 30624 14176
rect 30560 14116 30564 14172
rect 30564 14116 30620 14172
rect 30620 14116 30624 14172
rect 30560 14112 30624 14116
rect 30640 14172 30704 14176
rect 30640 14116 30644 14172
rect 30644 14116 30700 14172
rect 30700 14116 30704 14172
rect 30640 14112 30704 14116
rect 59848 14172 59912 14176
rect 59848 14116 59852 14172
rect 59852 14116 59908 14172
rect 59908 14116 59912 14172
rect 59848 14112 59912 14116
rect 59928 14172 59992 14176
rect 59928 14116 59932 14172
rect 59932 14116 59988 14172
rect 59988 14116 59992 14172
rect 59928 14112 59992 14116
rect 60008 14172 60072 14176
rect 60008 14116 60012 14172
rect 60012 14116 60068 14172
rect 60068 14116 60072 14172
rect 60008 14112 60072 14116
rect 60088 14172 60152 14176
rect 60088 14116 60092 14172
rect 60092 14116 60148 14172
rect 60148 14116 60152 14172
rect 60088 14112 60152 14116
rect 89296 14172 89360 14176
rect 89296 14116 89300 14172
rect 89300 14116 89356 14172
rect 89356 14116 89360 14172
rect 89296 14112 89360 14116
rect 89376 14172 89440 14176
rect 89376 14116 89380 14172
rect 89380 14116 89436 14172
rect 89436 14116 89440 14172
rect 89376 14112 89440 14116
rect 89456 14172 89520 14176
rect 89456 14116 89460 14172
rect 89460 14116 89516 14172
rect 89516 14116 89520 14172
rect 89456 14112 89520 14116
rect 89536 14172 89600 14176
rect 89536 14116 89540 14172
rect 89540 14116 89596 14172
rect 89596 14116 89600 14172
rect 89536 14112 89600 14116
rect 15676 13628 15740 13632
rect 15676 13572 15680 13628
rect 15680 13572 15736 13628
rect 15736 13572 15740 13628
rect 15676 13568 15740 13572
rect 15756 13628 15820 13632
rect 15756 13572 15760 13628
rect 15760 13572 15816 13628
rect 15816 13572 15820 13628
rect 15756 13568 15820 13572
rect 15836 13628 15900 13632
rect 15836 13572 15840 13628
rect 15840 13572 15896 13628
rect 15896 13572 15900 13628
rect 15836 13568 15900 13572
rect 15916 13628 15980 13632
rect 15916 13572 15920 13628
rect 15920 13572 15976 13628
rect 15976 13572 15980 13628
rect 15916 13568 15980 13572
rect 45124 13628 45188 13632
rect 45124 13572 45128 13628
rect 45128 13572 45184 13628
rect 45184 13572 45188 13628
rect 45124 13568 45188 13572
rect 45204 13628 45268 13632
rect 45204 13572 45208 13628
rect 45208 13572 45264 13628
rect 45264 13572 45268 13628
rect 45204 13568 45268 13572
rect 45284 13628 45348 13632
rect 45284 13572 45288 13628
rect 45288 13572 45344 13628
rect 45344 13572 45348 13628
rect 45284 13568 45348 13572
rect 45364 13628 45428 13632
rect 45364 13572 45368 13628
rect 45368 13572 45424 13628
rect 45424 13572 45428 13628
rect 45364 13568 45428 13572
rect 74572 13628 74636 13632
rect 74572 13572 74576 13628
rect 74576 13572 74632 13628
rect 74632 13572 74636 13628
rect 74572 13568 74636 13572
rect 74652 13628 74716 13632
rect 74652 13572 74656 13628
rect 74656 13572 74712 13628
rect 74712 13572 74716 13628
rect 74652 13568 74716 13572
rect 74732 13628 74796 13632
rect 74732 13572 74736 13628
rect 74736 13572 74792 13628
rect 74792 13572 74796 13628
rect 74732 13568 74796 13572
rect 74812 13628 74876 13632
rect 74812 13572 74816 13628
rect 74816 13572 74872 13628
rect 74872 13572 74876 13628
rect 74812 13568 74876 13572
rect 104020 13628 104084 13632
rect 104020 13572 104024 13628
rect 104024 13572 104080 13628
rect 104080 13572 104084 13628
rect 104020 13568 104084 13572
rect 104100 13628 104164 13632
rect 104100 13572 104104 13628
rect 104104 13572 104160 13628
rect 104160 13572 104164 13628
rect 104100 13568 104164 13572
rect 104180 13628 104244 13632
rect 104180 13572 104184 13628
rect 104184 13572 104240 13628
rect 104240 13572 104244 13628
rect 104180 13568 104244 13572
rect 104260 13628 104324 13632
rect 104260 13572 104264 13628
rect 104264 13572 104320 13628
rect 104320 13572 104324 13628
rect 104260 13568 104324 13572
rect 30400 13084 30464 13088
rect 30400 13028 30404 13084
rect 30404 13028 30460 13084
rect 30460 13028 30464 13084
rect 30400 13024 30464 13028
rect 30480 13084 30544 13088
rect 30480 13028 30484 13084
rect 30484 13028 30540 13084
rect 30540 13028 30544 13084
rect 30480 13024 30544 13028
rect 30560 13084 30624 13088
rect 30560 13028 30564 13084
rect 30564 13028 30620 13084
rect 30620 13028 30624 13084
rect 30560 13024 30624 13028
rect 30640 13084 30704 13088
rect 30640 13028 30644 13084
rect 30644 13028 30700 13084
rect 30700 13028 30704 13084
rect 30640 13024 30704 13028
rect 59848 13084 59912 13088
rect 59848 13028 59852 13084
rect 59852 13028 59908 13084
rect 59908 13028 59912 13084
rect 59848 13024 59912 13028
rect 59928 13084 59992 13088
rect 59928 13028 59932 13084
rect 59932 13028 59988 13084
rect 59988 13028 59992 13084
rect 59928 13024 59992 13028
rect 60008 13084 60072 13088
rect 60008 13028 60012 13084
rect 60012 13028 60068 13084
rect 60068 13028 60072 13084
rect 60008 13024 60072 13028
rect 60088 13084 60152 13088
rect 60088 13028 60092 13084
rect 60092 13028 60148 13084
rect 60148 13028 60152 13084
rect 60088 13024 60152 13028
rect 89296 13084 89360 13088
rect 89296 13028 89300 13084
rect 89300 13028 89356 13084
rect 89356 13028 89360 13084
rect 89296 13024 89360 13028
rect 89376 13084 89440 13088
rect 89376 13028 89380 13084
rect 89380 13028 89436 13084
rect 89436 13028 89440 13084
rect 89376 13024 89440 13028
rect 89456 13084 89520 13088
rect 89456 13028 89460 13084
rect 89460 13028 89516 13084
rect 89516 13028 89520 13084
rect 89456 13024 89520 13028
rect 89536 13084 89600 13088
rect 89536 13028 89540 13084
rect 89540 13028 89596 13084
rect 89596 13028 89600 13084
rect 89536 13024 89600 13028
rect 15676 12540 15740 12544
rect 15676 12484 15680 12540
rect 15680 12484 15736 12540
rect 15736 12484 15740 12540
rect 15676 12480 15740 12484
rect 15756 12540 15820 12544
rect 15756 12484 15760 12540
rect 15760 12484 15816 12540
rect 15816 12484 15820 12540
rect 15756 12480 15820 12484
rect 15836 12540 15900 12544
rect 15836 12484 15840 12540
rect 15840 12484 15896 12540
rect 15896 12484 15900 12540
rect 15836 12480 15900 12484
rect 15916 12540 15980 12544
rect 15916 12484 15920 12540
rect 15920 12484 15976 12540
rect 15976 12484 15980 12540
rect 15916 12480 15980 12484
rect 45124 12540 45188 12544
rect 45124 12484 45128 12540
rect 45128 12484 45184 12540
rect 45184 12484 45188 12540
rect 45124 12480 45188 12484
rect 45204 12540 45268 12544
rect 45204 12484 45208 12540
rect 45208 12484 45264 12540
rect 45264 12484 45268 12540
rect 45204 12480 45268 12484
rect 45284 12540 45348 12544
rect 45284 12484 45288 12540
rect 45288 12484 45344 12540
rect 45344 12484 45348 12540
rect 45284 12480 45348 12484
rect 45364 12540 45428 12544
rect 45364 12484 45368 12540
rect 45368 12484 45424 12540
rect 45424 12484 45428 12540
rect 45364 12480 45428 12484
rect 74572 12540 74636 12544
rect 74572 12484 74576 12540
rect 74576 12484 74632 12540
rect 74632 12484 74636 12540
rect 74572 12480 74636 12484
rect 74652 12540 74716 12544
rect 74652 12484 74656 12540
rect 74656 12484 74712 12540
rect 74712 12484 74716 12540
rect 74652 12480 74716 12484
rect 74732 12540 74796 12544
rect 74732 12484 74736 12540
rect 74736 12484 74792 12540
rect 74792 12484 74796 12540
rect 74732 12480 74796 12484
rect 74812 12540 74876 12544
rect 74812 12484 74816 12540
rect 74816 12484 74872 12540
rect 74872 12484 74876 12540
rect 74812 12480 74876 12484
rect 104020 12540 104084 12544
rect 104020 12484 104024 12540
rect 104024 12484 104080 12540
rect 104080 12484 104084 12540
rect 104020 12480 104084 12484
rect 104100 12540 104164 12544
rect 104100 12484 104104 12540
rect 104104 12484 104160 12540
rect 104160 12484 104164 12540
rect 104100 12480 104164 12484
rect 104180 12540 104244 12544
rect 104180 12484 104184 12540
rect 104184 12484 104240 12540
rect 104240 12484 104244 12540
rect 104180 12480 104244 12484
rect 104260 12540 104324 12544
rect 104260 12484 104264 12540
rect 104264 12484 104320 12540
rect 104320 12484 104324 12540
rect 104260 12480 104324 12484
rect 30400 11996 30464 12000
rect 30400 11940 30404 11996
rect 30404 11940 30460 11996
rect 30460 11940 30464 11996
rect 30400 11936 30464 11940
rect 30480 11996 30544 12000
rect 30480 11940 30484 11996
rect 30484 11940 30540 11996
rect 30540 11940 30544 11996
rect 30480 11936 30544 11940
rect 30560 11996 30624 12000
rect 30560 11940 30564 11996
rect 30564 11940 30620 11996
rect 30620 11940 30624 11996
rect 30560 11936 30624 11940
rect 30640 11996 30704 12000
rect 30640 11940 30644 11996
rect 30644 11940 30700 11996
rect 30700 11940 30704 11996
rect 30640 11936 30704 11940
rect 59848 11996 59912 12000
rect 59848 11940 59852 11996
rect 59852 11940 59908 11996
rect 59908 11940 59912 11996
rect 59848 11936 59912 11940
rect 59928 11996 59992 12000
rect 59928 11940 59932 11996
rect 59932 11940 59988 11996
rect 59988 11940 59992 11996
rect 59928 11936 59992 11940
rect 60008 11996 60072 12000
rect 60008 11940 60012 11996
rect 60012 11940 60068 11996
rect 60068 11940 60072 11996
rect 60008 11936 60072 11940
rect 60088 11996 60152 12000
rect 60088 11940 60092 11996
rect 60092 11940 60148 11996
rect 60148 11940 60152 11996
rect 60088 11936 60152 11940
rect 89296 11996 89360 12000
rect 89296 11940 89300 11996
rect 89300 11940 89356 11996
rect 89356 11940 89360 11996
rect 89296 11936 89360 11940
rect 89376 11996 89440 12000
rect 89376 11940 89380 11996
rect 89380 11940 89436 11996
rect 89436 11940 89440 11996
rect 89376 11936 89440 11940
rect 89456 11996 89520 12000
rect 89456 11940 89460 11996
rect 89460 11940 89516 11996
rect 89516 11940 89520 11996
rect 89456 11936 89520 11940
rect 89536 11996 89600 12000
rect 89536 11940 89540 11996
rect 89540 11940 89596 11996
rect 89596 11940 89600 11996
rect 89536 11936 89600 11940
rect 15676 11452 15740 11456
rect 15676 11396 15680 11452
rect 15680 11396 15736 11452
rect 15736 11396 15740 11452
rect 15676 11392 15740 11396
rect 15756 11452 15820 11456
rect 15756 11396 15760 11452
rect 15760 11396 15816 11452
rect 15816 11396 15820 11452
rect 15756 11392 15820 11396
rect 15836 11452 15900 11456
rect 15836 11396 15840 11452
rect 15840 11396 15896 11452
rect 15896 11396 15900 11452
rect 15836 11392 15900 11396
rect 15916 11452 15980 11456
rect 15916 11396 15920 11452
rect 15920 11396 15976 11452
rect 15976 11396 15980 11452
rect 15916 11392 15980 11396
rect 45124 11452 45188 11456
rect 45124 11396 45128 11452
rect 45128 11396 45184 11452
rect 45184 11396 45188 11452
rect 45124 11392 45188 11396
rect 45204 11452 45268 11456
rect 45204 11396 45208 11452
rect 45208 11396 45264 11452
rect 45264 11396 45268 11452
rect 45204 11392 45268 11396
rect 45284 11452 45348 11456
rect 45284 11396 45288 11452
rect 45288 11396 45344 11452
rect 45344 11396 45348 11452
rect 45284 11392 45348 11396
rect 45364 11452 45428 11456
rect 45364 11396 45368 11452
rect 45368 11396 45424 11452
rect 45424 11396 45428 11452
rect 45364 11392 45428 11396
rect 74572 11452 74636 11456
rect 74572 11396 74576 11452
rect 74576 11396 74632 11452
rect 74632 11396 74636 11452
rect 74572 11392 74636 11396
rect 74652 11452 74716 11456
rect 74652 11396 74656 11452
rect 74656 11396 74712 11452
rect 74712 11396 74716 11452
rect 74652 11392 74716 11396
rect 74732 11452 74796 11456
rect 74732 11396 74736 11452
rect 74736 11396 74792 11452
rect 74792 11396 74796 11452
rect 74732 11392 74796 11396
rect 74812 11452 74876 11456
rect 74812 11396 74816 11452
rect 74816 11396 74872 11452
rect 74872 11396 74876 11452
rect 74812 11392 74876 11396
rect 104020 11452 104084 11456
rect 104020 11396 104024 11452
rect 104024 11396 104080 11452
rect 104080 11396 104084 11452
rect 104020 11392 104084 11396
rect 104100 11452 104164 11456
rect 104100 11396 104104 11452
rect 104104 11396 104160 11452
rect 104160 11396 104164 11452
rect 104100 11392 104164 11396
rect 104180 11452 104244 11456
rect 104180 11396 104184 11452
rect 104184 11396 104240 11452
rect 104240 11396 104244 11452
rect 104180 11392 104244 11396
rect 104260 11452 104324 11456
rect 104260 11396 104264 11452
rect 104264 11396 104320 11452
rect 104320 11396 104324 11452
rect 104260 11392 104324 11396
rect 30400 10908 30464 10912
rect 30400 10852 30404 10908
rect 30404 10852 30460 10908
rect 30460 10852 30464 10908
rect 30400 10848 30464 10852
rect 30480 10908 30544 10912
rect 30480 10852 30484 10908
rect 30484 10852 30540 10908
rect 30540 10852 30544 10908
rect 30480 10848 30544 10852
rect 30560 10908 30624 10912
rect 30560 10852 30564 10908
rect 30564 10852 30620 10908
rect 30620 10852 30624 10908
rect 30560 10848 30624 10852
rect 30640 10908 30704 10912
rect 30640 10852 30644 10908
rect 30644 10852 30700 10908
rect 30700 10852 30704 10908
rect 30640 10848 30704 10852
rect 59848 10908 59912 10912
rect 59848 10852 59852 10908
rect 59852 10852 59908 10908
rect 59908 10852 59912 10908
rect 59848 10848 59912 10852
rect 59928 10908 59992 10912
rect 59928 10852 59932 10908
rect 59932 10852 59988 10908
rect 59988 10852 59992 10908
rect 59928 10848 59992 10852
rect 60008 10908 60072 10912
rect 60008 10852 60012 10908
rect 60012 10852 60068 10908
rect 60068 10852 60072 10908
rect 60008 10848 60072 10852
rect 60088 10908 60152 10912
rect 60088 10852 60092 10908
rect 60092 10852 60148 10908
rect 60148 10852 60152 10908
rect 60088 10848 60152 10852
rect 89296 10908 89360 10912
rect 89296 10852 89300 10908
rect 89300 10852 89356 10908
rect 89356 10852 89360 10908
rect 89296 10848 89360 10852
rect 89376 10908 89440 10912
rect 89376 10852 89380 10908
rect 89380 10852 89436 10908
rect 89436 10852 89440 10908
rect 89376 10848 89440 10852
rect 89456 10908 89520 10912
rect 89456 10852 89460 10908
rect 89460 10852 89516 10908
rect 89516 10852 89520 10908
rect 89456 10848 89520 10852
rect 89536 10908 89600 10912
rect 89536 10852 89540 10908
rect 89540 10852 89596 10908
rect 89596 10852 89600 10908
rect 89536 10848 89600 10852
rect 15676 10364 15740 10368
rect 15676 10308 15680 10364
rect 15680 10308 15736 10364
rect 15736 10308 15740 10364
rect 15676 10304 15740 10308
rect 15756 10364 15820 10368
rect 15756 10308 15760 10364
rect 15760 10308 15816 10364
rect 15816 10308 15820 10364
rect 15756 10304 15820 10308
rect 15836 10364 15900 10368
rect 15836 10308 15840 10364
rect 15840 10308 15896 10364
rect 15896 10308 15900 10364
rect 15836 10304 15900 10308
rect 15916 10364 15980 10368
rect 15916 10308 15920 10364
rect 15920 10308 15976 10364
rect 15976 10308 15980 10364
rect 15916 10304 15980 10308
rect 45124 10364 45188 10368
rect 45124 10308 45128 10364
rect 45128 10308 45184 10364
rect 45184 10308 45188 10364
rect 45124 10304 45188 10308
rect 45204 10364 45268 10368
rect 45204 10308 45208 10364
rect 45208 10308 45264 10364
rect 45264 10308 45268 10364
rect 45204 10304 45268 10308
rect 45284 10364 45348 10368
rect 45284 10308 45288 10364
rect 45288 10308 45344 10364
rect 45344 10308 45348 10364
rect 45284 10304 45348 10308
rect 45364 10364 45428 10368
rect 45364 10308 45368 10364
rect 45368 10308 45424 10364
rect 45424 10308 45428 10364
rect 45364 10304 45428 10308
rect 74572 10364 74636 10368
rect 74572 10308 74576 10364
rect 74576 10308 74632 10364
rect 74632 10308 74636 10364
rect 74572 10304 74636 10308
rect 74652 10364 74716 10368
rect 74652 10308 74656 10364
rect 74656 10308 74712 10364
rect 74712 10308 74716 10364
rect 74652 10304 74716 10308
rect 74732 10364 74796 10368
rect 74732 10308 74736 10364
rect 74736 10308 74792 10364
rect 74792 10308 74796 10364
rect 74732 10304 74796 10308
rect 74812 10364 74876 10368
rect 74812 10308 74816 10364
rect 74816 10308 74872 10364
rect 74872 10308 74876 10364
rect 74812 10304 74876 10308
rect 104020 10364 104084 10368
rect 104020 10308 104024 10364
rect 104024 10308 104080 10364
rect 104080 10308 104084 10364
rect 104020 10304 104084 10308
rect 104100 10364 104164 10368
rect 104100 10308 104104 10364
rect 104104 10308 104160 10364
rect 104160 10308 104164 10364
rect 104100 10304 104164 10308
rect 104180 10364 104244 10368
rect 104180 10308 104184 10364
rect 104184 10308 104240 10364
rect 104240 10308 104244 10364
rect 104180 10304 104244 10308
rect 104260 10364 104324 10368
rect 104260 10308 104264 10364
rect 104264 10308 104320 10364
rect 104320 10308 104324 10364
rect 104260 10304 104324 10308
rect 30400 9820 30464 9824
rect 30400 9764 30404 9820
rect 30404 9764 30460 9820
rect 30460 9764 30464 9820
rect 30400 9760 30464 9764
rect 30480 9820 30544 9824
rect 30480 9764 30484 9820
rect 30484 9764 30540 9820
rect 30540 9764 30544 9820
rect 30480 9760 30544 9764
rect 30560 9820 30624 9824
rect 30560 9764 30564 9820
rect 30564 9764 30620 9820
rect 30620 9764 30624 9820
rect 30560 9760 30624 9764
rect 30640 9820 30704 9824
rect 30640 9764 30644 9820
rect 30644 9764 30700 9820
rect 30700 9764 30704 9820
rect 30640 9760 30704 9764
rect 59848 9820 59912 9824
rect 59848 9764 59852 9820
rect 59852 9764 59908 9820
rect 59908 9764 59912 9820
rect 59848 9760 59912 9764
rect 59928 9820 59992 9824
rect 59928 9764 59932 9820
rect 59932 9764 59988 9820
rect 59988 9764 59992 9820
rect 59928 9760 59992 9764
rect 60008 9820 60072 9824
rect 60008 9764 60012 9820
rect 60012 9764 60068 9820
rect 60068 9764 60072 9820
rect 60008 9760 60072 9764
rect 60088 9820 60152 9824
rect 60088 9764 60092 9820
rect 60092 9764 60148 9820
rect 60148 9764 60152 9820
rect 60088 9760 60152 9764
rect 89296 9820 89360 9824
rect 89296 9764 89300 9820
rect 89300 9764 89356 9820
rect 89356 9764 89360 9820
rect 89296 9760 89360 9764
rect 89376 9820 89440 9824
rect 89376 9764 89380 9820
rect 89380 9764 89436 9820
rect 89436 9764 89440 9820
rect 89376 9760 89440 9764
rect 89456 9820 89520 9824
rect 89456 9764 89460 9820
rect 89460 9764 89516 9820
rect 89516 9764 89520 9820
rect 89456 9760 89520 9764
rect 89536 9820 89600 9824
rect 89536 9764 89540 9820
rect 89540 9764 89596 9820
rect 89596 9764 89600 9820
rect 89536 9760 89600 9764
rect 15676 9276 15740 9280
rect 15676 9220 15680 9276
rect 15680 9220 15736 9276
rect 15736 9220 15740 9276
rect 15676 9216 15740 9220
rect 15756 9276 15820 9280
rect 15756 9220 15760 9276
rect 15760 9220 15816 9276
rect 15816 9220 15820 9276
rect 15756 9216 15820 9220
rect 15836 9276 15900 9280
rect 15836 9220 15840 9276
rect 15840 9220 15896 9276
rect 15896 9220 15900 9276
rect 15836 9216 15900 9220
rect 15916 9276 15980 9280
rect 15916 9220 15920 9276
rect 15920 9220 15976 9276
rect 15976 9220 15980 9276
rect 15916 9216 15980 9220
rect 45124 9276 45188 9280
rect 45124 9220 45128 9276
rect 45128 9220 45184 9276
rect 45184 9220 45188 9276
rect 45124 9216 45188 9220
rect 45204 9276 45268 9280
rect 45204 9220 45208 9276
rect 45208 9220 45264 9276
rect 45264 9220 45268 9276
rect 45204 9216 45268 9220
rect 45284 9276 45348 9280
rect 45284 9220 45288 9276
rect 45288 9220 45344 9276
rect 45344 9220 45348 9276
rect 45284 9216 45348 9220
rect 45364 9276 45428 9280
rect 45364 9220 45368 9276
rect 45368 9220 45424 9276
rect 45424 9220 45428 9276
rect 45364 9216 45428 9220
rect 74572 9276 74636 9280
rect 74572 9220 74576 9276
rect 74576 9220 74632 9276
rect 74632 9220 74636 9276
rect 74572 9216 74636 9220
rect 74652 9276 74716 9280
rect 74652 9220 74656 9276
rect 74656 9220 74712 9276
rect 74712 9220 74716 9276
rect 74652 9216 74716 9220
rect 74732 9276 74796 9280
rect 74732 9220 74736 9276
rect 74736 9220 74792 9276
rect 74792 9220 74796 9276
rect 74732 9216 74796 9220
rect 74812 9276 74876 9280
rect 74812 9220 74816 9276
rect 74816 9220 74872 9276
rect 74872 9220 74876 9276
rect 74812 9216 74876 9220
rect 104020 9276 104084 9280
rect 104020 9220 104024 9276
rect 104024 9220 104080 9276
rect 104080 9220 104084 9276
rect 104020 9216 104084 9220
rect 104100 9276 104164 9280
rect 104100 9220 104104 9276
rect 104104 9220 104160 9276
rect 104160 9220 104164 9276
rect 104100 9216 104164 9220
rect 104180 9276 104244 9280
rect 104180 9220 104184 9276
rect 104184 9220 104240 9276
rect 104240 9220 104244 9276
rect 104180 9216 104244 9220
rect 104260 9276 104324 9280
rect 104260 9220 104264 9276
rect 104264 9220 104320 9276
rect 104320 9220 104324 9276
rect 104260 9216 104324 9220
rect 30400 8732 30464 8736
rect 30400 8676 30404 8732
rect 30404 8676 30460 8732
rect 30460 8676 30464 8732
rect 30400 8672 30464 8676
rect 30480 8732 30544 8736
rect 30480 8676 30484 8732
rect 30484 8676 30540 8732
rect 30540 8676 30544 8732
rect 30480 8672 30544 8676
rect 30560 8732 30624 8736
rect 30560 8676 30564 8732
rect 30564 8676 30620 8732
rect 30620 8676 30624 8732
rect 30560 8672 30624 8676
rect 30640 8732 30704 8736
rect 30640 8676 30644 8732
rect 30644 8676 30700 8732
rect 30700 8676 30704 8732
rect 30640 8672 30704 8676
rect 59848 8732 59912 8736
rect 59848 8676 59852 8732
rect 59852 8676 59908 8732
rect 59908 8676 59912 8732
rect 59848 8672 59912 8676
rect 59928 8732 59992 8736
rect 59928 8676 59932 8732
rect 59932 8676 59988 8732
rect 59988 8676 59992 8732
rect 59928 8672 59992 8676
rect 60008 8732 60072 8736
rect 60008 8676 60012 8732
rect 60012 8676 60068 8732
rect 60068 8676 60072 8732
rect 60008 8672 60072 8676
rect 60088 8732 60152 8736
rect 60088 8676 60092 8732
rect 60092 8676 60148 8732
rect 60148 8676 60152 8732
rect 60088 8672 60152 8676
rect 89296 8732 89360 8736
rect 89296 8676 89300 8732
rect 89300 8676 89356 8732
rect 89356 8676 89360 8732
rect 89296 8672 89360 8676
rect 89376 8732 89440 8736
rect 89376 8676 89380 8732
rect 89380 8676 89436 8732
rect 89436 8676 89440 8732
rect 89376 8672 89440 8676
rect 89456 8732 89520 8736
rect 89456 8676 89460 8732
rect 89460 8676 89516 8732
rect 89516 8676 89520 8732
rect 89456 8672 89520 8676
rect 89536 8732 89600 8736
rect 89536 8676 89540 8732
rect 89540 8676 89596 8732
rect 89596 8676 89600 8732
rect 89536 8672 89600 8676
rect 15676 8188 15740 8192
rect 15676 8132 15680 8188
rect 15680 8132 15736 8188
rect 15736 8132 15740 8188
rect 15676 8128 15740 8132
rect 15756 8188 15820 8192
rect 15756 8132 15760 8188
rect 15760 8132 15816 8188
rect 15816 8132 15820 8188
rect 15756 8128 15820 8132
rect 15836 8188 15900 8192
rect 15836 8132 15840 8188
rect 15840 8132 15896 8188
rect 15896 8132 15900 8188
rect 15836 8128 15900 8132
rect 15916 8188 15980 8192
rect 15916 8132 15920 8188
rect 15920 8132 15976 8188
rect 15976 8132 15980 8188
rect 15916 8128 15980 8132
rect 45124 8188 45188 8192
rect 45124 8132 45128 8188
rect 45128 8132 45184 8188
rect 45184 8132 45188 8188
rect 45124 8128 45188 8132
rect 45204 8188 45268 8192
rect 45204 8132 45208 8188
rect 45208 8132 45264 8188
rect 45264 8132 45268 8188
rect 45204 8128 45268 8132
rect 45284 8188 45348 8192
rect 45284 8132 45288 8188
rect 45288 8132 45344 8188
rect 45344 8132 45348 8188
rect 45284 8128 45348 8132
rect 45364 8188 45428 8192
rect 45364 8132 45368 8188
rect 45368 8132 45424 8188
rect 45424 8132 45428 8188
rect 45364 8128 45428 8132
rect 74572 8188 74636 8192
rect 74572 8132 74576 8188
rect 74576 8132 74632 8188
rect 74632 8132 74636 8188
rect 74572 8128 74636 8132
rect 74652 8188 74716 8192
rect 74652 8132 74656 8188
rect 74656 8132 74712 8188
rect 74712 8132 74716 8188
rect 74652 8128 74716 8132
rect 74732 8188 74796 8192
rect 74732 8132 74736 8188
rect 74736 8132 74792 8188
rect 74792 8132 74796 8188
rect 74732 8128 74796 8132
rect 74812 8188 74876 8192
rect 74812 8132 74816 8188
rect 74816 8132 74872 8188
rect 74872 8132 74876 8188
rect 74812 8128 74876 8132
rect 104020 8188 104084 8192
rect 104020 8132 104024 8188
rect 104024 8132 104080 8188
rect 104080 8132 104084 8188
rect 104020 8128 104084 8132
rect 104100 8188 104164 8192
rect 104100 8132 104104 8188
rect 104104 8132 104160 8188
rect 104160 8132 104164 8188
rect 104100 8128 104164 8132
rect 104180 8188 104244 8192
rect 104180 8132 104184 8188
rect 104184 8132 104240 8188
rect 104240 8132 104244 8188
rect 104180 8128 104244 8132
rect 104260 8188 104324 8192
rect 104260 8132 104264 8188
rect 104264 8132 104320 8188
rect 104320 8132 104324 8188
rect 104260 8128 104324 8132
rect 30400 7644 30464 7648
rect 30400 7588 30404 7644
rect 30404 7588 30460 7644
rect 30460 7588 30464 7644
rect 30400 7584 30464 7588
rect 30480 7644 30544 7648
rect 30480 7588 30484 7644
rect 30484 7588 30540 7644
rect 30540 7588 30544 7644
rect 30480 7584 30544 7588
rect 30560 7644 30624 7648
rect 30560 7588 30564 7644
rect 30564 7588 30620 7644
rect 30620 7588 30624 7644
rect 30560 7584 30624 7588
rect 30640 7644 30704 7648
rect 30640 7588 30644 7644
rect 30644 7588 30700 7644
rect 30700 7588 30704 7644
rect 30640 7584 30704 7588
rect 59848 7644 59912 7648
rect 59848 7588 59852 7644
rect 59852 7588 59908 7644
rect 59908 7588 59912 7644
rect 59848 7584 59912 7588
rect 59928 7644 59992 7648
rect 59928 7588 59932 7644
rect 59932 7588 59988 7644
rect 59988 7588 59992 7644
rect 59928 7584 59992 7588
rect 60008 7644 60072 7648
rect 60008 7588 60012 7644
rect 60012 7588 60068 7644
rect 60068 7588 60072 7644
rect 60008 7584 60072 7588
rect 60088 7644 60152 7648
rect 60088 7588 60092 7644
rect 60092 7588 60148 7644
rect 60148 7588 60152 7644
rect 60088 7584 60152 7588
rect 89296 7644 89360 7648
rect 89296 7588 89300 7644
rect 89300 7588 89356 7644
rect 89356 7588 89360 7644
rect 89296 7584 89360 7588
rect 89376 7644 89440 7648
rect 89376 7588 89380 7644
rect 89380 7588 89436 7644
rect 89436 7588 89440 7644
rect 89376 7584 89440 7588
rect 89456 7644 89520 7648
rect 89456 7588 89460 7644
rect 89460 7588 89516 7644
rect 89516 7588 89520 7644
rect 89456 7584 89520 7588
rect 89536 7644 89600 7648
rect 89536 7588 89540 7644
rect 89540 7588 89596 7644
rect 89596 7588 89600 7644
rect 89536 7584 89600 7588
rect 15676 7100 15740 7104
rect 15676 7044 15680 7100
rect 15680 7044 15736 7100
rect 15736 7044 15740 7100
rect 15676 7040 15740 7044
rect 15756 7100 15820 7104
rect 15756 7044 15760 7100
rect 15760 7044 15816 7100
rect 15816 7044 15820 7100
rect 15756 7040 15820 7044
rect 15836 7100 15900 7104
rect 15836 7044 15840 7100
rect 15840 7044 15896 7100
rect 15896 7044 15900 7100
rect 15836 7040 15900 7044
rect 15916 7100 15980 7104
rect 15916 7044 15920 7100
rect 15920 7044 15976 7100
rect 15976 7044 15980 7100
rect 15916 7040 15980 7044
rect 45124 7100 45188 7104
rect 45124 7044 45128 7100
rect 45128 7044 45184 7100
rect 45184 7044 45188 7100
rect 45124 7040 45188 7044
rect 45204 7100 45268 7104
rect 45204 7044 45208 7100
rect 45208 7044 45264 7100
rect 45264 7044 45268 7100
rect 45204 7040 45268 7044
rect 45284 7100 45348 7104
rect 45284 7044 45288 7100
rect 45288 7044 45344 7100
rect 45344 7044 45348 7100
rect 45284 7040 45348 7044
rect 45364 7100 45428 7104
rect 45364 7044 45368 7100
rect 45368 7044 45424 7100
rect 45424 7044 45428 7100
rect 45364 7040 45428 7044
rect 74572 7100 74636 7104
rect 74572 7044 74576 7100
rect 74576 7044 74632 7100
rect 74632 7044 74636 7100
rect 74572 7040 74636 7044
rect 74652 7100 74716 7104
rect 74652 7044 74656 7100
rect 74656 7044 74712 7100
rect 74712 7044 74716 7100
rect 74652 7040 74716 7044
rect 74732 7100 74796 7104
rect 74732 7044 74736 7100
rect 74736 7044 74792 7100
rect 74792 7044 74796 7100
rect 74732 7040 74796 7044
rect 74812 7100 74876 7104
rect 74812 7044 74816 7100
rect 74816 7044 74872 7100
rect 74872 7044 74876 7100
rect 74812 7040 74876 7044
rect 104020 7100 104084 7104
rect 104020 7044 104024 7100
rect 104024 7044 104080 7100
rect 104080 7044 104084 7100
rect 104020 7040 104084 7044
rect 104100 7100 104164 7104
rect 104100 7044 104104 7100
rect 104104 7044 104160 7100
rect 104160 7044 104164 7100
rect 104100 7040 104164 7044
rect 104180 7100 104244 7104
rect 104180 7044 104184 7100
rect 104184 7044 104240 7100
rect 104240 7044 104244 7100
rect 104180 7040 104244 7044
rect 104260 7100 104324 7104
rect 104260 7044 104264 7100
rect 104264 7044 104320 7100
rect 104320 7044 104324 7100
rect 104260 7040 104324 7044
rect 30400 6556 30464 6560
rect 30400 6500 30404 6556
rect 30404 6500 30460 6556
rect 30460 6500 30464 6556
rect 30400 6496 30464 6500
rect 30480 6556 30544 6560
rect 30480 6500 30484 6556
rect 30484 6500 30540 6556
rect 30540 6500 30544 6556
rect 30480 6496 30544 6500
rect 30560 6556 30624 6560
rect 30560 6500 30564 6556
rect 30564 6500 30620 6556
rect 30620 6500 30624 6556
rect 30560 6496 30624 6500
rect 30640 6556 30704 6560
rect 30640 6500 30644 6556
rect 30644 6500 30700 6556
rect 30700 6500 30704 6556
rect 30640 6496 30704 6500
rect 59848 6556 59912 6560
rect 59848 6500 59852 6556
rect 59852 6500 59908 6556
rect 59908 6500 59912 6556
rect 59848 6496 59912 6500
rect 59928 6556 59992 6560
rect 59928 6500 59932 6556
rect 59932 6500 59988 6556
rect 59988 6500 59992 6556
rect 59928 6496 59992 6500
rect 60008 6556 60072 6560
rect 60008 6500 60012 6556
rect 60012 6500 60068 6556
rect 60068 6500 60072 6556
rect 60008 6496 60072 6500
rect 60088 6556 60152 6560
rect 60088 6500 60092 6556
rect 60092 6500 60148 6556
rect 60148 6500 60152 6556
rect 60088 6496 60152 6500
rect 89296 6556 89360 6560
rect 89296 6500 89300 6556
rect 89300 6500 89356 6556
rect 89356 6500 89360 6556
rect 89296 6496 89360 6500
rect 89376 6556 89440 6560
rect 89376 6500 89380 6556
rect 89380 6500 89436 6556
rect 89436 6500 89440 6556
rect 89376 6496 89440 6500
rect 89456 6556 89520 6560
rect 89456 6500 89460 6556
rect 89460 6500 89516 6556
rect 89516 6500 89520 6556
rect 89456 6496 89520 6500
rect 89536 6556 89600 6560
rect 89536 6500 89540 6556
rect 89540 6500 89596 6556
rect 89596 6500 89600 6556
rect 89536 6496 89600 6500
rect 15676 6012 15740 6016
rect 15676 5956 15680 6012
rect 15680 5956 15736 6012
rect 15736 5956 15740 6012
rect 15676 5952 15740 5956
rect 15756 6012 15820 6016
rect 15756 5956 15760 6012
rect 15760 5956 15816 6012
rect 15816 5956 15820 6012
rect 15756 5952 15820 5956
rect 15836 6012 15900 6016
rect 15836 5956 15840 6012
rect 15840 5956 15896 6012
rect 15896 5956 15900 6012
rect 15836 5952 15900 5956
rect 15916 6012 15980 6016
rect 15916 5956 15920 6012
rect 15920 5956 15976 6012
rect 15976 5956 15980 6012
rect 15916 5952 15980 5956
rect 45124 6012 45188 6016
rect 45124 5956 45128 6012
rect 45128 5956 45184 6012
rect 45184 5956 45188 6012
rect 45124 5952 45188 5956
rect 45204 6012 45268 6016
rect 45204 5956 45208 6012
rect 45208 5956 45264 6012
rect 45264 5956 45268 6012
rect 45204 5952 45268 5956
rect 45284 6012 45348 6016
rect 45284 5956 45288 6012
rect 45288 5956 45344 6012
rect 45344 5956 45348 6012
rect 45284 5952 45348 5956
rect 45364 6012 45428 6016
rect 45364 5956 45368 6012
rect 45368 5956 45424 6012
rect 45424 5956 45428 6012
rect 45364 5952 45428 5956
rect 74572 6012 74636 6016
rect 74572 5956 74576 6012
rect 74576 5956 74632 6012
rect 74632 5956 74636 6012
rect 74572 5952 74636 5956
rect 74652 6012 74716 6016
rect 74652 5956 74656 6012
rect 74656 5956 74712 6012
rect 74712 5956 74716 6012
rect 74652 5952 74716 5956
rect 74732 6012 74796 6016
rect 74732 5956 74736 6012
rect 74736 5956 74792 6012
rect 74792 5956 74796 6012
rect 74732 5952 74796 5956
rect 74812 6012 74876 6016
rect 74812 5956 74816 6012
rect 74816 5956 74872 6012
rect 74872 5956 74876 6012
rect 74812 5952 74876 5956
rect 104020 6012 104084 6016
rect 104020 5956 104024 6012
rect 104024 5956 104080 6012
rect 104080 5956 104084 6012
rect 104020 5952 104084 5956
rect 104100 6012 104164 6016
rect 104100 5956 104104 6012
rect 104104 5956 104160 6012
rect 104160 5956 104164 6012
rect 104100 5952 104164 5956
rect 104180 6012 104244 6016
rect 104180 5956 104184 6012
rect 104184 5956 104240 6012
rect 104240 5956 104244 6012
rect 104180 5952 104244 5956
rect 104260 6012 104324 6016
rect 104260 5956 104264 6012
rect 104264 5956 104320 6012
rect 104320 5956 104324 6012
rect 104260 5952 104324 5956
rect 30400 5468 30464 5472
rect 30400 5412 30404 5468
rect 30404 5412 30460 5468
rect 30460 5412 30464 5468
rect 30400 5408 30464 5412
rect 30480 5468 30544 5472
rect 30480 5412 30484 5468
rect 30484 5412 30540 5468
rect 30540 5412 30544 5468
rect 30480 5408 30544 5412
rect 30560 5468 30624 5472
rect 30560 5412 30564 5468
rect 30564 5412 30620 5468
rect 30620 5412 30624 5468
rect 30560 5408 30624 5412
rect 30640 5468 30704 5472
rect 30640 5412 30644 5468
rect 30644 5412 30700 5468
rect 30700 5412 30704 5468
rect 30640 5408 30704 5412
rect 59848 5468 59912 5472
rect 59848 5412 59852 5468
rect 59852 5412 59908 5468
rect 59908 5412 59912 5468
rect 59848 5408 59912 5412
rect 59928 5468 59992 5472
rect 59928 5412 59932 5468
rect 59932 5412 59988 5468
rect 59988 5412 59992 5468
rect 59928 5408 59992 5412
rect 60008 5468 60072 5472
rect 60008 5412 60012 5468
rect 60012 5412 60068 5468
rect 60068 5412 60072 5468
rect 60008 5408 60072 5412
rect 60088 5468 60152 5472
rect 60088 5412 60092 5468
rect 60092 5412 60148 5468
rect 60148 5412 60152 5468
rect 60088 5408 60152 5412
rect 89296 5468 89360 5472
rect 89296 5412 89300 5468
rect 89300 5412 89356 5468
rect 89356 5412 89360 5468
rect 89296 5408 89360 5412
rect 89376 5468 89440 5472
rect 89376 5412 89380 5468
rect 89380 5412 89436 5468
rect 89436 5412 89440 5468
rect 89376 5408 89440 5412
rect 89456 5468 89520 5472
rect 89456 5412 89460 5468
rect 89460 5412 89516 5468
rect 89516 5412 89520 5468
rect 89456 5408 89520 5412
rect 89536 5468 89600 5472
rect 89536 5412 89540 5468
rect 89540 5412 89596 5468
rect 89596 5412 89600 5468
rect 89536 5408 89600 5412
rect 15676 4924 15740 4928
rect 15676 4868 15680 4924
rect 15680 4868 15736 4924
rect 15736 4868 15740 4924
rect 15676 4864 15740 4868
rect 15756 4924 15820 4928
rect 15756 4868 15760 4924
rect 15760 4868 15816 4924
rect 15816 4868 15820 4924
rect 15756 4864 15820 4868
rect 15836 4924 15900 4928
rect 15836 4868 15840 4924
rect 15840 4868 15896 4924
rect 15896 4868 15900 4924
rect 15836 4864 15900 4868
rect 15916 4924 15980 4928
rect 15916 4868 15920 4924
rect 15920 4868 15976 4924
rect 15976 4868 15980 4924
rect 15916 4864 15980 4868
rect 45124 4924 45188 4928
rect 45124 4868 45128 4924
rect 45128 4868 45184 4924
rect 45184 4868 45188 4924
rect 45124 4864 45188 4868
rect 45204 4924 45268 4928
rect 45204 4868 45208 4924
rect 45208 4868 45264 4924
rect 45264 4868 45268 4924
rect 45204 4864 45268 4868
rect 45284 4924 45348 4928
rect 45284 4868 45288 4924
rect 45288 4868 45344 4924
rect 45344 4868 45348 4924
rect 45284 4864 45348 4868
rect 45364 4924 45428 4928
rect 45364 4868 45368 4924
rect 45368 4868 45424 4924
rect 45424 4868 45428 4924
rect 45364 4864 45428 4868
rect 74572 4924 74636 4928
rect 74572 4868 74576 4924
rect 74576 4868 74632 4924
rect 74632 4868 74636 4924
rect 74572 4864 74636 4868
rect 74652 4924 74716 4928
rect 74652 4868 74656 4924
rect 74656 4868 74712 4924
rect 74712 4868 74716 4924
rect 74652 4864 74716 4868
rect 74732 4924 74796 4928
rect 74732 4868 74736 4924
rect 74736 4868 74792 4924
rect 74792 4868 74796 4924
rect 74732 4864 74796 4868
rect 74812 4924 74876 4928
rect 74812 4868 74816 4924
rect 74816 4868 74872 4924
rect 74872 4868 74876 4924
rect 74812 4864 74876 4868
rect 104020 4924 104084 4928
rect 104020 4868 104024 4924
rect 104024 4868 104080 4924
rect 104080 4868 104084 4924
rect 104020 4864 104084 4868
rect 104100 4924 104164 4928
rect 104100 4868 104104 4924
rect 104104 4868 104160 4924
rect 104160 4868 104164 4924
rect 104100 4864 104164 4868
rect 104180 4924 104244 4928
rect 104180 4868 104184 4924
rect 104184 4868 104240 4924
rect 104240 4868 104244 4924
rect 104180 4864 104244 4868
rect 104260 4924 104324 4928
rect 104260 4868 104264 4924
rect 104264 4868 104320 4924
rect 104320 4868 104324 4924
rect 104260 4864 104324 4868
rect 30400 4380 30464 4384
rect 30400 4324 30404 4380
rect 30404 4324 30460 4380
rect 30460 4324 30464 4380
rect 30400 4320 30464 4324
rect 30480 4380 30544 4384
rect 30480 4324 30484 4380
rect 30484 4324 30540 4380
rect 30540 4324 30544 4380
rect 30480 4320 30544 4324
rect 30560 4380 30624 4384
rect 30560 4324 30564 4380
rect 30564 4324 30620 4380
rect 30620 4324 30624 4380
rect 30560 4320 30624 4324
rect 30640 4380 30704 4384
rect 30640 4324 30644 4380
rect 30644 4324 30700 4380
rect 30700 4324 30704 4380
rect 30640 4320 30704 4324
rect 59848 4380 59912 4384
rect 59848 4324 59852 4380
rect 59852 4324 59908 4380
rect 59908 4324 59912 4380
rect 59848 4320 59912 4324
rect 59928 4380 59992 4384
rect 59928 4324 59932 4380
rect 59932 4324 59988 4380
rect 59988 4324 59992 4380
rect 59928 4320 59992 4324
rect 60008 4380 60072 4384
rect 60008 4324 60012 4380
rect 60012 4324 60068 4380
rect 60068 4324 60072 4380
rect 60008 4320 60072 4324
rect 60088 4380 60152 4384
rect 60088 4324 60092 4380
rect 60092 4324 60148 4380
rect 60148 4324 60152 4380
rect 60088 4320 60152 4324
rect 89296 4380 89360 4384
rect 89296 4324 89300 4380
rect 89300 4324 89356 4380
rect 89356 4324 89360 4380
rect 89296 4320 89360 4324
rect 89376 4380 89440 4384
rect 89376 4324 89380 4380
rect 89380 4324 89436 4380
rect 89436 4324 89440 4380
rect 89376 4320 89440 4324
rect 89456 4380 89520 4384
rect 89456 4324 89460 4380
rect 89460 4324 89516 4380
rect 89516 4324 89520 4380
rect 89456 4320 89520 4324
rect 89536 4380 89600 4384
rect 89536 4324 89540 4380
rect 89540 4324 89596 4380
rect 89596 4324 89600 4380
rect 89536 4320 89600 4324
rect 15676 3836 15740 3840
rect 15676 3780 15680 3836
rect 15680 3780 15736 3836
rect 15736 3780 15740 3836
rect 15676 3776 15740 3780
rect 15756 3836 15820 3840
rect 15756 3780 15760 3836
rect 15760 3780 15816 3836
rect 15816 3780 15820 3836
rect 15756 3776 15820 3780
rect 15836 3836 15900 3840
rect 15836 3780 15840 3836
rect 15840 3780 15896 3836
rect 15896 3780 15900 3836
rect 15836 3776 15900 3780
rect 15916 3836 15980 3840
rect 15916 3780 15920 3836
rect 15920 3780 15976 3836
rect 15976 3780 15980 3836
rect 15916 3776 15980 3780
rect 45124 3836 45188 3840
rect 45124 3780 45128 3836
rect 45128 3780 45184 3836
rect 45184 3780 45188 3836
rect 45124 3776 45188 3780
rect 45204 3836 45268 3840
rect 45204 3780 45208 3836
rect 45208 3780 45264 3836
rect 45264 3780 45268 3836
rect 45204 3776 45268 3780
rect 45284 3836 45348 3840
rect 45284 3780 45288 3836
rect 45288 3780 45344 3836
rect 45344 3780 45348 3836
rect 45284 3776 45348 3780
rect 45364 3836 45428 3840
rect 45364 3780 45368 3836
rect 45368 3780 45424 3836
rect 45424 3780 45428 3836
rect 45364 3776 45428 3780
rect 74572 3836 74636 3840
rect 74572 3780 74576 3836
rect 74576 3780 74632 3836
rect 74632 3780 74636 3836
rect 74572 3776 74636 3780
rect 74652 3836 74716 3840
rect 74652 3780 74656 3836
rect 74656 3780 74712 3836
rect 74712 3780 74716 3836
rect 74652 3776 74716 3780
rect 74732 3836 74796 3840
rect 74732 3780 74736 3836
rect 74736 3780 74792 3836
rect 74792 3780 74796 3836
rect 74732 3776 74796 3780
rect 74812 3836 74876 3840
rect 74812 3780 74816 3836
rect 74816 3780 74872 3836
rect 74872 3780 74876 3836
rect 74812 3776 74876 3780
rect 104020 3836 104084 3840
rect 104020 3780 104024 3836
rect 104024 3780 104080 3836
rect 104080 3780 104084 3836
rect 104020 3776 104084 3780
rect 104100 3836 104164 3840
rect 104100 3780 104104 3836
rect 104104 3780 104160 3836
rect 104160 3780 104164 3836
rect 104100 3776 104164 3780
rect 104180 3836 104244 3840
rect 104180 3780 104184 3836
rect 104184 3780 104240 3836
rect 104240 3780 104244 3836
rect 104180 3776 104244 3780
rect 104260 3836 104324 3840
rect 104260 3780 104264 3836
rect 104264 3780 104320 3836
rect 104320 3780 104324 3836
rect 104260 3776 104324 3780
rect 30400 3292 30464 3296
rect 30400 3236 30404 3292
rect 30404 3236 30460 3292
rect 30460 3236 30464 3292
rect 30400 3232 30464 3236
rect 30480 3292 30544 3296
rect 30480 3236 30484 3292
rect 30484 3236 30540 3292
rect 30540 3236 30544 3292
rect 30480 3232 30544 3236
rect 30560 3292 30624 3296
rect 30560 3236 30564 3292
rect 30564 3236 30620 3292
rect 30620 3236 30624 3292
rect 30560 3232 30624 3236
rect 30640 3292 30704 3296
rect 30640 3236 30644 3292
rect 30644 3236 30700 3292
rect 30700 3236 30704 3292
rect 30640 3232 30704 3236
rect 59848 3292 59912 3296
rect 59848 3236 59852 3292
rect 59852 3236 59908 3292
rect 59908 3236 59912 3292
rect 59848 3232 59912 3236
rect 59928 3292 59992 3296
rect 59928 3236 59932 3292
rect 59932 3236 59988 3292
rect 59988 3236 59992 3292
rect 59928 3232 59992 3236
rect 60008 3292 60072 3296
rect 60008 3236 60012 3292
rect 60012 3236 60068 3292
rect 60068 3236 60072 3292
rect 60008 3232 60072 3236
rect 60088 3292 60152 3296
rect 60088 3236 60092 3292
rect 60092 3236 60148 3292
rect 60148 3236 60152 3292
rect 60088 3232 60152 3236
rect 89296 3292 89360 3296
rect 89296 3236 89300 3292
rect 89300 3236 89356 3292
rect 89356 3236 89360 3292
rect 89296 3232 89360 3236
rect 89376 3292 89440 3296
rect 89376 3236 89380 3292
rect 89380 3236 89436 3292
rect 89436 3236 89440 3292
rect 89376 3232 89440 3236
rect 89456 3292 89520 3296
rect 89456 3236 89460 3292
rect 89460 3236 89516 3292
rect 89516 3236 89520 3292
rect 89456 3232 89520 3236
rect 89536 3292 89600 3296
rect 89536 3236 89540 3292
rect 89540 3236 89596 3292
rect 89596 3236 89600 3292
rect 89536 3232 89600 3236
rect 15676 2748 15740 2752
rect 15676 2692 15680 2748
rect 15680 2692 15736 2748
rect 15736 2692 15740 2748
rect 15676 2688 15740 2692
rect 15756 2748 15820 2752
rect 15756 2692 15760 2748
rect 15760 2692 15816 2748
rect 15816 2692 15820 2748
rect 15756 2688 15820 2692
rect 15836 2748 15900 2752
rect 15836 2692 15840 2748
rect 15840 2692 15896 2748
rect 15896 2692 15900 2748
rect 15836 2688 15900 2692
rect 15916 2748 15980 2752
rect 15916 2692 15920 2748
rect 15920 2692 15976 2748
rect 15976 2692 15980 2748
rect 15916 2688 15980 2692
rect 45124 2748 45188 2752
rect 45124 2692 45128 2748
rect 45128 2692 45184 2748
rect 45184 2692 45188 2748
rect 45124 2688 45188 2692
rect 45204 2748 45268 2752
rect 45204 2692 45208 2748
rect 45208 2692 45264 2748
rect 45264 2692 45268 2748
rect 45204 2688 45268 2692
rect 45284 2748 45348 2752
rect 45284 2692 45288 2748
rect 45288 2692 45344 2748
rect 45344 2692 45348 2748
rect 45284 2688 45348 2692
rect 45364 2748 45428 2752
rect 45364 2692 45368 2748
rect 45368 2692 45424 2748
rect 45424 2692 45428 2748
rect 45364 2688 45428 2692
rect 74572 2748 74636 2752
rect 74572 2692 74576 2748
rect 74576 2692 74632 2748
rect 74632 2692 74636 2748
rect 74572 2688 74636 2692
rect 74652 2748 74716 2752
rect 74652 2692 74656 2748
rect 74656 2692 74712 2748
rect 74712 2692 74716 2748
rect 74652 2688 74716 2692
rect 74732 2748 74796 2752
rect 74732 2692 74736 2748
rect 74736 2692 74792 2748
rect 74792 2692 74796 2748
rect 74732 2688 74796 2692
rect 74812 2748 74876 2752
rect 74812 2692 74816 2748
rect 74816 2692 74872 2748
rect 74872 2692 74876 2748
rect 74812 2688 74876 2692
rect 104020 2748 104084 2752
rect 104020 2692 104024 2748
rect 104024 2692 104080 2748
rect 104080 2692 104084 2748
rect 104020 2688 104084 2692
rect 104100 2748 104164 2752
rect 104100 2692 104104 2748
rect 104104 2692 104160 2748
rect 104160 2692 104164 2748
rect 104100 2688 104164 2692
rect 104180 2748 104244 2752
rect 104180 2692 104184 2748
rect 104184 2692 104240 2748
rect 104240 2692 104244 2748
rect 104180 2688 104244 2692
rect 104260 2748 104324 2752
rect 104260 2692 104264 2748
rect 104264 2692 104320 2748
rect 104320 2692 104324 2748
rect 104260 2688 104324 2692
rect 30400 2204 30464 2208
rect 30400 2148 30404 2204
rect 30404 2148 30460 2204
rect 30460 2148 30464 2204
rect 30400 2144 30464 2148
rect 30480 2204 30544 2208
rect 30480 2148 30484 2204
rect 30484 2148 30540 2204
rect 30540 2148 30544 2204
rect 30480 2144 30544 2148
rect 30560 2204 30624 2208
rect 30560 2148 30564 2204
rect 30564 2148 30620 2204
rect 30620 2148 30624 2204
rect 30560 2144 30624 2148
rect 30640 2204 30704 2208
rect 30640 2148 30644 2204
rect 30644 2148 30700 2204
rect 30700 2148 30704 2204
rect 30640 2144 30704 2148
rect 59848 2204 59912 2208
rect 59848 2148 59852 2204
rect 59852 2148 59908 2204
rect 59908 2148 59912 2204
rect 59848 2144 59912 2148
rect 59928 2204 59992 2208
rect 59928 2148 59932 2204
rect 59932 2148 59988 2204
rect 59988 2148 59992 2204
rect 59928 2144 59992 2148
rect 60008 2204 60072 2208
rect 60008 2148 60012 2204
rect 60012 2148 60068 2204
rect 60068 2148 60072 2204
rect 60008 2144 60072 2148
rect 60088 2204 60152 2208
rect 60088 2148 60092 2204
rect 60092 2148 60148 2204
rect 60148 2148 60152 2204
rect 60088 2144 60152 2148
rect 89296 2204 89360 2208
rect 89296 2148 89300 2204
rect 89300 2148 89356 2204
rect 89356 2148 89360 2204
rect 89296 2144 89360 2148
rect 89376 2204 89440 2208
rect 89376 2148 89380 2204
rect 89380 2148 89436 2204
rect 89436 2148 89440 2204
rect 89376 2144 89440 2148
rect 89456 2204 89520 2208
rect 89456 2148 89460 2204
rect 89460 2148 89516 2204
rect 89516 2148 89520 2204
rect 89456 2144 89520 2148
rect 89536 2204 89600 2208
rect 89536 2148 89540 2204
rect 89540 2148 89596 2204
rect 89596 2148 89600 2204
rect 89536 2144 89600 2148
<< metal4 >>
rect 15668 27776 15988 27792
rect 15668 27712 15676 27776
rect 15740 27712 15756 27776
rect 15820 27712 15836 27776
rect 15900 27712 15916 27776
rect 15980 27712 15988 27776
rect 15668 26688 15988 27712
rect 15668 26624 15676 26688
rect 15740 26624 15756 26688
rect 15820 26624 15836 26688
rect 15900 26624 15916 26688
rect 15980 26624 15988 26688
rect 15668 25600 15988 26624
rect 15668 25536 15676 25600
rect 15740 25536 15756 25600
rect 15820 25536 15836 25600
rect 15900 25536 15916 25600
rect 15980 25536 15988 25600
rect 15668 24512 15988 25536
rect 15668 24448 15676 24512
rect 15740 24448 15756 24512
rect 15820 24448 15836 24512
rect 15900 24448 15916 24512
rect 15980 24448 15988 24512
rect 15668 23424 15988 24448
rect 15668 23360 15676 23424
rect 15740 23360 15756 23424
rect 15820 23360 15836 23424
rect 15900 23360 15916 23424
rect 15980 23360 15988 23424
rect 15668 22336 15988 23360
rect 15668 22272 15676 22336
rect 15740 22272 15756 22336
rect 15820 22272 15836 22336
rect 15900 22272 15916 22336
rect 15980 22272 15988 22336
rect 15668 21248 15988 22272
rect 15668 21184 15676 21248
rect 15740 21184 15756 21248
rect 15820 21184 15836 21248
rect 15900 21184 15916 21248
rect 15980 21184 15988 21248
rect 15668 20160 15988 21184
rect 15668 20096 15676 20160
rect 15740 20096 15756 20160
rect 15820 20096 15836 20160
rect 15900 20096 15916 20160
rect 15980 20096 15988 20160
rect 15668 19072 15988 20096
rect 15668 19008 15676 19072
rect 15740 19008 15756 19072
rect 15820 19008 15836 19072
rect 15900 19008 15916 19072
rect 15980 19008 15988 19072
rect 15668 17984 15988 19008
rect 15668 17920 15676 17984
rect 15740 17920 15756 17984
rect 15820 17920 15836 17984
rect 15900 17920 15916 17984
rect 15980 17920 15988 17984
rect 15668 16896 15988 17920
rect 15668 16832 15676 16896
rect 15740 16832 15756 16896
rect 15820 16832 15836 16896
rect 15900 16832 15916 16896
rect 15980 16832 15988 16896
rect 15668 15808 15988 16832
rect 15668 15744 15676 15808
rect 15740 15744 15756 15808
rect 15820 15744 15836 15808
rect 15900 15744 15916 15808
rect 15980 15744 15988 15808
rect 15668 14720 15988 15744
rect 15668 14656 15676 14720
rect 15740 14656 15756 14720
rect 15820 14656 15836 14720
rect 15900 14656 15916 14720
rect 15980 14656 15988 14720
rect 15668 13632 15988 14656
rect 15668 13568 15676 13632
rect 15740 13568 15756 13632
rect 15820 13568 15836 13632
rect 15900 13568 15916 13632
rect 15980 13568 15988 13632
rect 15668 12544 15988 13568
rect 15668 12480 15676 12544
rect 15740 12480 15756 12544
rect 15820 12480 15836 12544
rect 15900 12480 15916 12544
rect 15980 12480 15988 12544
rect 15668 11456 15988 12480
rect 15668 11392 15676 11456
rect 15740 11392 15756 11456
rect 15820 11392 15836 11456
rect 15900 11392 15916 11456
rect 15980 11392 15988 11456
rect 15668 10368 15988 11392
rect 15668 10304 15676 10368
rect 15740 10304 15756 10368
rect 15820 10304 15836 10368
rect 15900 10304 15916 10368
rect 15980 10304 15988 10368
rect 15668 9280 15988 10304
rect 15668 9216 15676 9280
rect 15740 9216 15756 9280
rect 15820 9216 15836 9280
rect 15900 9216 15916 9280
rect 15980 9216 15988 9280
rect 15668 8192 15988 9216
rect 15668 8128 15676 8192
rect 15740 8128 15756 8192
rect 15820 8128 15836 8192
rect 15900 8128 15916 8192
rect 15980 8128 15988 8192
rect 15668 7104 15988 8128
rect 15668 7040 15676 7104
rect 15740 7040 15756 7104
rect 15820 7040 15836 7104
rect 15900 7040 15916 7104
rect 15980 7040 15988 7104
rect 15668 6016 15988 7040
rect 15668 5952 15676 6016
rect 15740 5952 15756 6016
rect 15820 5952 15836 6016
rect 15900 5952 15916 6016
rect 15980 5952 15988 6016
rect 15668 4928 15988 5952
rect 15668 4864 15676 4928
rect 15740 4864 15756 4928
rect 15820 4864 15836 4928
rect 15900 4864 15916 4928
rect 15980 4864 15988 4928
rect 15668 3840 15988 4864
rect 15668 3776 15676 3840
rect 15740 3776 15756 3840
rect 15820 3776 15836 3840
rect 15900 3776 15916 3840
rect 15980 3776 15988 3840
rect 15668 2752 15988 3776
rect 15668 2688 15676 2752
rect 15740 2688 15756 2752
rect 15820 2688 15836 2752
rect 15900 2688 15916 2752
rect 15980 2688 15988 2752
rect 15668 2128 15988 2688
rect 30392 27232 30712 27792
rect 30392 27168 30400 27232
rect 30464 27168 30480 27232
rect 30544 27168 30560 27232
rect 30624 27168 30640 27232
rect 30704 27168 30712 27232
rect 30392 26144 30712 27168
rect 30392 26080 30400 26144
rect 30464 26080 30480 26144
rect 30544 26080 30560 26144
rect 30624 26080 30640 26144
rect 30704 26080 30712 26144
rect 30392 25056 30712 26080
rect 30392 24992 30400 25056
rect 30464 24992 30480 25056
rect 30544 24992 30560 25056
rect 30624 24992 30640 25056
rect 30704 24992 30712 25056
rect 30392 23968 30712 24992
rect 30392 23904 30400 23968
rect 30464 23904 30480 23968
rect 30544 23904 30560 23968
rect 30624 23904 30640 23968
rect 30704 23904 30712 23968
rect 30392 22880 30712 23904
rect 30392 22816 30400 22880
rect 30464 22816 30480 22880
rect 30544 22816 30560 22880
rect 30624 22816 30640 22880
rect 30704 22816 30712 22880
rect 30392 21792 30712 22816
rect 30392 21728 30400 21792
rect 30464 21728 30480 21792
rect 30544 21728 30560 21792
rect 30624 21728 30640 21792
rect 30704 21728 30712 21792
rect 30392 20704 30712 21728
rect 30392 20640 30400 20704
rect 30464 20640 30480 20704
rect 30544 20640 30560 20704
rect 30624 20640 30640 20704
rect 30704 20640 30712 20704
rect 30392 19616 30712 20640
rect 30392 19552 30400 19616
rect 30464 19552 30480 19616
rect 30544 19552 30560 19616
rect 30624 19552 30640 19616
rect 30704 19552 30712 19616
rect 30392 18528 30712 19552
rect 30392 18464 30400 18528
rect 30464 18464 30480 18528
rect 30544 18464 30560 18528
rect 30624 18464 30640 18528
rect 30704 18464 30712 18528
rect 30392 17440 30712 18464
rect 30392 17376 30400 17440
rect 30464 17376 30480 17440
rect 30544 17376 30560 17440
rect 30624 17376 30640 17440
rect 30704 17376 30712 17440
rect 30392 16352 30712 17376
rect 30392 16288 30400 16352
rect 30464 16288 30480 16352
rect 30544 16288 30560 16352
rect 30624 16288 30640 16352
rect 30704 16288 30712 16352
rect 30392 15264 30712 16288
rect 30392 15200 30400 15264
rect 30464 15200 30480 15264
rect 30544 15200 30560 15264
rect 30624 15200 30640 15264
rect 30704 15200 30712 15264
rect 30392 14176 30712 15200
rect 30392 14112 30400 14176
rect 30464 14112 30480 14176
rect 30544 14112 30560 14176
rect 30624 14112 30640 14176
rect 30704 14112 30712 14176
rect 30392 13088 30712 14112
rect 30392 13024 30400 13088
rect 30464 13024 30480 13088
rect 30544 13024 30560 13088
rect 30624 13024 30640 13088
rect 30704 13024 30712 13088
rect 30392 12000 30712 13024
rect 30392 11936 30400 12000
rect 30464 11936 30480 12000
rect 30544 11936 30560 12000
rect 30624 11936 30640 12000
rect 30704 11936 30712 12000
rect 30392 10912 30712 11936
rect 30392 10848 30400 10912
rect 30464 10848 30480 10912
rect 30544 10848 30560 10912
rect 30624 10848 30640 10912
rect 30704 10848 30712 10912
rect 30392 9824 30712 10848
rect 30392 9760 30400 9824
rect 30464 9760 30480 9824
rect 30544 9760 30560 9824
rect 30624 9760 30640 9824
rect 30704 9760 30712 9824
rect 30392 8736 30712 9760
rect 30392 8672 30400 8736
rect 30464 8672 30480 8736
rect 30544 8672 30560 8736
rect 30624 8672 30640 8736
rect 30704 8672 30712 8736
rect 30392 7648 30712 8672
rect 30392 7584 30400 7648
rect 30464 7584 30480 7648
rect 30544 7584 30560 7648
rect 30624 7584 30640 7648
rect 30704 7584 30712 7648
rect 30392 6560 30712 7584
rect 30392 6496 30400 6560
rect 30464 6496 30480 6560
rect 30544 6496 30560 6560
rect 30624 6496 30640 6560
rect 30704 6496 30712 6560
rect 30392 5472 30712 6496
rect 30392 5408 30400 5472
rect 30464 5408 30480 5472
rect 30544 5408 30560 5472
rect 30624 5408 30640 5472
rect 30704 5408 30712 5472
rect 30392 4384 30712 5408
rect 30392 4320 30400 4384
rect 30464 4320 30480 4384
rect 30544 4320 30560 4384
rect 30624 4320 30640 4384
rect 30704 4320 30712 4384
rect 30392 3296 30712 4320
rect 30392 3232 30400 3296
rect 30464 3232 30480 3296
rect 30544 3232 30560 3296
rect 30624 3232 30640 3296
rect 30704 3232 30712 3296
rect 30392 2208 30712 3232
rect 30392 2144 30400 2208
rect 30464 2144 30480 2208
rect 30544 2144 30560 2208
rect 30624 2144 30640 2208
rect 30704 2144 30712 2208
rect 30392 2128 30712 2144
rect 45116 27776 45436 27792
rect 45116 27712 45124 27776
rect 45188 27712 45204 27776
rect 45268 27712 45284 27776
rect 45348 27712 45364 27776
rect 45428 27712 45436 27776
rect 45116 26688 45436 27712
rect 45116 26624 45124 26688
rect 45188 26624 45204 26688
rect 45268 26624 45284 26688
rect 45348 26624 45364 26688
rect 45428 26624 45436 26688
rect 45116 25600 45436 26624
rect 45116 25536 45124 25600
rect 45188 25536 45204 25600
rect 45268 25536 45284 25600
rect 45348 25536 45364 25600
rect 45428 25536 45436 25600
rect 45116 24512 45436 25536
rect 45116 24448 45124 24512
rect 45188 24448 45204 24512
rect 45268 24448 45284 24512
rect 45348 24448 45364 24512
rect 45428 24448 45436 24512
rect 45116 23424 45436 24448
rect 45116 23360 45124 23424
rect 45188 23360 45204 23424
rect 45268 23360 45284 23424
rect 45348 23360 45364 23424
rect 45428 23360 45436 23424
rect 45116 22336 45436 23360
rect 45116 22272 45124 22336
rect 45188 22272 45204 22336
rect 45268 22272 45284 22336
rect 45348 22272 45364 22336
rect 45428 22272 45436 22336
rect 45116 21248 45436 22272
rect 45116 21184 45124 21248
rect 45188 21184 45204 21248
rect 45268 21184 45284 21248
rect 45348 21184 45364 21248
rect 45428 21184 45436 21248
rect 45116 20160 45436 21184
rect 45116 20096 45124 20160
rect 45188 20096 45204 20160
rect 45268 20096 45284 20160
rect 45348 20096 45364 20160
rect 45428 20096 45436 20160
rect 45116 19072 45436 20096
rect 45116 19008 45124 19072
rect 45188 19008 45204 19072
rect 45268 19008 45284 19072
rect 45348 19008 45364 19072
rect 45428 19008 45436 19072
rect 45116 17984 45436 19008
rect 45116 17920 45124 17984
rect 45188 17920 45204 17984
rect 45268 17920 45284 17984
rect 45348 17920 45364 17984
rect 45428 17920 45436 17984
rect 45116 16896 45436 17920
rect 45116 16832 45124 16896
rect 45188 16832 45204 16896
rect 45268 16832 45284 16896
rect 45348 16832 45364 16896
rect 45428 16832 45436 16896
rect 45116 15808 45436 16832
rect 45116 15744 45124 15808
rect 45188 15744 45204 15808
rect 45268 15744 45284 15808
rect 45348 15744 45364 15808
rect 45428 15744 45436 15808
rect 45116 14720 45436 15744
rect 45116 14656 45124 14720
rect 45188 14656 45204 14720
rect 45268 14656 45284 14720
rect 45348 14656 45364 14720
rect 45428 14656 45436 14720
rect 45116 13632 45436 14656
rect 45116 13568 45124 13632
rect 45188 13568 45204 13632
rect 45268 13568 45284 13632
rect 45348 13568 45364 13632
rect 45428 13568 45436 13632
rect 45116 12544 45436 13568
rect 45116 12480 45124 12544
rect 45188 12480 45204 12544
rect 45268 12480 45284 12544
rect 45348 12480 45364 12544
rect 45428 12480 45436 12544
rect 45116 11456 45436 12480
rect 45116 11392 45124 11456
rect 45188 11392 45204 11456
rect 45268 11392 45284 11456
rect 45348 11392 45364 11456
rect 45428 11392 45436 11456
rect 45116 10368 45436 11392
rect 45116 10304 45124 10368
rect 45188 10304 45204 10368
rect 45268 10304 45284 10368
rect 45348 10304 45364 10368
rect 45428 10304 45436 10368
rect 45116 9280 45436 10304
rect 45116 9216 45124 9280
rect 45188 9216 45204 9280
rect 45268 9216 45284 9280
rect 45348 9216 45364 9280
rect 45428 9216 45436 9280
rect 45116 8192 45436 9216
rect 45116 8128 45124 8192
rect 45188 8128 45204 8192
rect 45268 8128 45284 8192
rect 45348 8128 45364 8192
rect 45428 8128 45436 8192
rect 45116 7104 45436 8128
rect 45116 7040 45124 7104
rect 45188 7040 45204 7104
rect 45268 7040 45284 7104
rect 45348 7040 45364 7104
rect 45428 7040 45436 7104
rect 45116 6016 45436 7040
rect 45116 5952 45124 6016
rect 45188 5952 45204 6016
rect 45268 5952 45284 6016
rect 45348 5952 45364 6016
rect 45428 5952 45436 6016
rect 45116 4928 45436 5952
rect 45116 4864 45124 4928
rect 45188 4864 45204 4928
rect 45268 4864 45284 4928
rect 45348 4864 45364 4928
rect 45428 4864 45436 4928
rect 45116 3840 45436 4864
rect 45116 3776 45124 3840
rect 45188 3776 45204 3840
rect 45268 3776 45284 3840
rect 45348 3776 45364 3840
rect 45428 3776 45436 3840
rect 45116 2752 45436 3776
rect 45116 2688 45124 2752
rect 45188 2688 45204 2752
rect 45268 2688 45284 2752
rect 45348 2688 45364 2752
rect 45428 2688 45436 2752
rect 45116 2128 45436 2688
rect 59840 27232 60160 27792
rect 59840 27168 59848 27232
rect 59912 27168 59928 27232
rect 59992 27168 60008 27232
rect 60072 27168 60088 27232
rect 60152 27168 60160 27232
rect 59840 26144 60160 27168
rect 74564 27776 74884 27792
rect 74564 27712 74572 27776
rect 74636 27712 74652 27776
rect 74716 27712 74732 27776
rect 74796 27712 74812 27776
rect 74876 27712 74884 27776
rect 70350 26830 70778 26890
rect 70350 26757 70410 26830
rect 70347 26756 70413 26757
rect 70347 26692 70348 26756
rect 70412 26692 70413 26756
rect 70347 26691 70413 26692
rect 70718 26349 70778 26830
rect 74564 26688 74884 27712
rect 74564 26624 74572 26688
rect 74636 26624 74652 26688
rect 74716 26624 74732 26688
rect 74796 26624 74812 26688
rect 74876 26624 74884 26688
rect 70715 26348 70781 26349
rect 70715 26284 70716 26348
rect 70780 26284 70781 26348
rect 70715 26283 70781 26284
rect 59840 26080 59848 26144
rect 59912 26080 59928 26144
rect 59992 26080 60008 26144
rect 60072 26080 60088 26144
rect 60152 26080 60160 26144
rect 59840 25056 60160 26080
rect 59840 24992 59848 25056
rect 59912 24992 59928 25056
rect 59992 24992 60008 25056
rect 60072 24992 60088 25056
rect 60152 24992 60160 25056
rect 59840 23968 60160 24992
rect 59840 23904 59848 23968
rect 59912 23904 59928 23968
rect 59992 23904 60008 23968
rect 60072 23904 60088 23968
rect 60152 23904 60160 23968
rect 59840 22880 60160 23904
rect 59840 22816 59848 22880
rect 59912 22816 59928 22880
rect 59992 22816 60008 22880
rect 60072 22816 60088 22880
rect 60152 22816 60160 22880
rect 59840 21792 60160 22816
rect 59840 21728 59848 21792
rect 59912 21728 59928 21792
rect 59992 21728 60008 21792
rect 60072 21728 60088 21792
rect 60152 21728 60160 21792
rect 59840 20704 60160 21728
rect 59840 20640 59848 20704
rect 59912 20640 59928 20704
rect 59992 20640 60008 20704
rect 60072 20640 60088 20704
rect 60152 20640 60160 20704
rect 59840 19616 60160 20640
rect 59840 19552 59848 19616
rect 59912 19552 59928 19616
rect 59992 19552 60008 19616
rect 60072 19552 60088 19616
rect 60152 19552 60160 19616
rect 59840 18528 60160 19552
rect 59840 18464 59848 18528
rect 59912 18464 59928 18528
rect 59992 18464 60008 18528
rect 60072 18464 60088 18528
rect 60152 18464 60160 18528
rect 59840 17440 60160 18464
rect 59840 17376 59848 17440
rect 59912 17376 59928 17440
rect 59992 17376 60008 17440
rect 60072 17376 60088 17440
rect 60152 17376 60160 17440
rect 59840 16352 60160 17376
rect 59840 16288 59848 16352
rect 59912 16288 59928 16352
rect 59992 16288 60008 16352
rect 60072 16288 60088 16352
rect 60152 16288 60160 16352
rect 59840 15264 60160 16288
rect 59840 15200 59848 15264
rect 59912 15200 59928 15264
rect 59992 15200 60008 15264
rect 60072 15200 60088 15264
rect 60152 15200 60160 15264
rect 59840 14176 60160 15200
rect 59840 14112 59848 14176
rect 59912 14112 59928 14176
rect 59992 14112 60008 14176
rect 60072 14112 60088 14176
rect 60152 14112 60160 14176
rect 59840 13088 60160 14112
rect 59840 13024 59848 13088
rect 59912 13024 59928 13088
rect 59992 13024 60008 13088
rect 60072 13024 60088 13088
rect 60152 13024 60160 13088
rect 59840 12000 60160 13024
rect 59840 11936 59848 12000
rect 59912 11936 59928 12000
rect 59992 11936 60008 12000
rect 60072 11936 60088 12000
rect 60152 11936 60160 12000
rect 59840 10912 60160 11936
rect 59840 10848 59848 10912
rect 59912 10848 59928 10912
rect 59992 10848 60008 10912
rect 60072 10848 60088 10912
rect 60152 10848 60160 10912
rect 59840 9824 60160 10848
rect 59840 9760 59848 9824
rect 59912 9760 59928 9824
rect 59992 9760 60008 9824
rect 60072 9760 60088 9824
rect 60152 9760 60160 9824
rect 59840 8736 60160 9760
rect 59840 8672 59848 8736
rect 59912 8672 59928 8736
rect 59992 8672 60008 8736
rect 60072 8672 60088 8736
rect 60152 8672 60160 8736
rect 59840 7648 60160 8672
rect 59840 7584 59848 7648
rect 59912 7584 59928 7648
rect 59992 7584 60008 7648
rect 60072 7584 60088 7648
rect 60152 7584 60160 7648
rect 59840 6560 60160 7584
rect 59840 6496 59848 6560
rect 59912 6496 59928 6560
rect 59992 6496 60008 6560
rect 60072 6496 60088 6560
rect 60152 6496 60160 6560
rect 59840 5472 60160 6496
rect 59840 5408 59848 5472
rect 59912 5408 59928 5472
rect 59992 5408 60008 5472
rect 60072 5408 60088 5472
rect 60152 5408 60160 5472
rect 59840 4384 60160 5408
rect 59840 4320 59848 4384
rect 59912 4320 59928 4384
rect 59992 4320 60008 4384
rect 60072 4320 60088 4384
rect 60152 4320 60160 4384
rect 59840 3296 60160 4320
rect 59840 3232 59848 3296
rect 59912 3232 59928 3296
rect 59992 3232 60008 3296
rect 60072 3232 60088 3296
rect 60152 3232 60160 3296
rect 59840 2208 60160 3232
rect 59840 2144 59848 2208
rect 59912 2144 59928 2208
rect 59992 2144 60008 2208
rect 60072 2144 60088 2208
rect 60152 2144 60160 2208
rect 59840 2128 60160 2144
rect 74564 25600 74884 26624
rect 74564 25536 74572 25600
rect 74636 25536 74652 25600
rect 74716 25536 74732 25600
rect 74796 25536 74812 25600
rect 74876 25536 74884 25600
rect 74564 24512 74884 25536
rect 74564 24448 74572 24512
rect 74636 24448 74652 24512
rect 74716 24448 74732 24512
rect 74796 24448 74812 24512
rect 74876 24448 74884 24512
rect 74564 23424 74884 24448
rect 74564 23360 74572 23424
rect 74636 23360 74652 23424
rect 74716 23360 74732 23424
rect 74796 23360 74812 23424
rect 74876 23360 74884 23424
rect 74564 22336 74884 23360
rect 74564 22272 74572 22336
rect 74636 22272 74652 22336
rect 74716 22272 74732 22336
rect 74796 22272 74812 22336
rect 74876 22272 74884 22336
rect 74564 21248 74884 22272
rect 74564 21184 74572 21248
rect 74636 21184 74652 21248
rect 74716 21184 74732 21248
rect 74796 21184 74812 21248
rect 74876 21184 74884 21248
rect 74564 20160 74884 21184
rect 74564 20096 74572 20160
rect 74636 20096 74652 20160
rect 74716 20096 74732 20160
rect 74796 20096 74812 20160
rect 74876 20096 74884 20160
rect 74564 19072 74884 20096
rect 74564 19008 74572 19072
rect 74636 19008 74652 19072
rect 74716 19008 74732 19072
rect 74796 19008 74812 19072
rect 74876 19008 74884 19072
rect 74564 17984 74884 19008
rect 74564 17920 74572 17984
rect 74636 17920 74652 17984
rect 74716 17920 74732 17984
rect 74796 17920 74812 17984
rect 74876 17920 74884 17984
rect 74564 16896 74884 17920
rect 74564 16832 74572 16896
rect 74636 16832 74652 16896
rect 74716 16832 74732 16896
rect 74796 16832 74812 16896
rect 74876 16832 74884 16896
rect 74564 15808 74884 16832
rect 74564 15744 74572 15808
rect 74636 15744 74652 15808
rect 74716 15744 74732 15808
rect 74796 15744 74812 15808
rect 74876 15744 74884 15808
rect 74564 14720 74884 15744
rect 74564 14656 74572 14720
rect 74636 14656 74652 14720
rect 74716 14656 74732 14720
rect 74796 14656 74812 14720
rect 74876 14656 74884 14720
rect 74564 13632 74884 14656
rect 74564 13568 74572 13632
rect 74636 13568 74652 13632
rect 74716 13568 74732 13632
rect 74796 13568 74812 13632
rect 74876 13568 74884 13632
rect 74564 12544 74884 13568
rect 74564 12480 74572 12544
rect 74636 12480 74652 12544
rect 74716 12480 74732 12544
rect 74796 12480 74812 12544
rect 74876 12480 74884 12544
rect 74564 11456 74884 12480
rect 74564 11392 74572 11456
rect 74636 11392 74652 11456
rect 74716 11392 74732 11456
rect 74796 11392 74812 11456
rect 74876 11392 74884 11456
rect 74564 10368 74884 11392
rect 74564 10304 74572 10368
rect 74636 10304 74652 10368
rect 74716 10304 74732 10368
rect 74796 10304 74812 10368
rect 74876 10304 74884 10368
rect 74564 9280 74884 10304
rect 74564 9216 74572 9280
rect 74636 9216 74652 9280
rect 74716 9216 74732 9280
rect 74796 9216 74812 9280
rect 74876 9216 74884 9280
rect 74564 8192 74884 9216
rect 74564 8128 74572 8192
rect 74636 8128 74652 8192
rect 74716 8128 74732 8192
rect 74796 8128 74812 8192
rect 74876 8128 74884 8192
rect 74564 7104 74884 8128
rect 74564 7040 74572 7104
rect 74636 7040 74652 7104
rect 74716 7040 74732 7104
rect 74796 7040 74812 7104
rect 74876 7040 74884 7104
rect 74564 6016 74884 7040
rect 74564 5952 74572 6016
rect 74636 5952 74652 6016
rect 74716 5952 74732 6016
rect 74796 5952 74812 6016
rect 74876 5952 74884 6016
rect 74564 4928 74884 5952
rect 74564 4864 74572 4928
rect 74636 4864 74652 4928
rect 74716 4864 74732 4928
rect 74796 4864 74812 4928
rect 74876 4864 74884 4928
rect 74564 3840 74884 4864
rect 74564 3776 74572 3840
rect 74636 3776 74652 3840
rect 74716 3776 74732 3840
rect 74796 3776 74812 3840
rect 74876 3776 74884 3840
rect 74564 2752 74884 3776
rect 74564 2688 74572 2752
rect 74636 2688 74652 2752
rect 74716 2688 74732 2752
rect 74796 2688 74812 2752
rect 74876 2688 74884 2752
rect 74564 2128 74884 2688
rect 89288 27232 89608 27792
rect 89288 27168 89296 27232
rect 89360 27168 89376 27232
rect 89440 27168 89456 27232
rect 89520 27168 89536 27232
rect 89600 27168 89608 27232
rect 89288 26144 89608 27168
rect 89288 26080 89296 26144
rect 89360 26080 89376 26144
rect 89440 26080 89456 26144
rect 89520 26080 89536 26144
rect 89600 26080 89608 26144
rect 89288 25056 89608 26080
rect 89288 24992 89296 25056
rect 89360 24992 89376 25056
rect 89440 24992 89456 25056
rect 89520 24992 89536 25056
rect 89600 24992 89608 25056
rect 89288 23968 89608 24992
rect 89288 23904 89296 23968
rect 89360 23904 89376 23968
rect 89440 23904 89456 23968
rect 89520 23904 89536 23968
rect 89600 23904 89608 23968
rect 89288 22880 89608 23904
rect 89288 22816 89296 22880
rect 89360 22816 89376 22880
rect 89440 22816 89456 22880
rect 89520 22816 89536 22880
rect 89600 22816 89608 22880
rect 89288 21792 89608 22816
rect 89288 21728 89296 21792
rect 89360 21728 89376 21792
rect 89440 21728 89456 21792
rect 89520 21728 89536 21792
rect 89600 21728 89608 21792
rect 89288 20704 89608 21728
rect 89288 20640 89296 20704
rect 89360 20640 89376 20704
rect 89440 20640 89456 20704
rect 89520 20640 89536 20704
rect 89600 20640 89608 20704
rect 89288 19616 89608 20640
rect 89288 19552 89296 19616
rect 89360 19552 89376 19616
rect 89440 19552 89456 19616
rect 89520 19552 89536 19616
rect 89600 19552 89608 19616
rect 89288 18528 89608 19552
rect 89288 18464 89296 18528
rect 89360 18464 89376 18528
rect 89440 18464 89456 18528
rect 89520 18464 89536 18528
rect 89600 18464 89608 18528
rect 89288 17440 89608 18464
rect 89288 17376 89296 17440
rect 89360 17376 89376 17440
rect 89440 17376 89456 17440
rect 89520 17376 89536 17440
rect 89600 17376 89608 17440
rect 89288 16352 89608 17376
rect 89288 16288 89296 16352
rect 89360 16288 89376 16352
rect 89440 16288 89456 16352
rect 89520 16288 89536 16352
rect 89600 16288 89608 16352
rect 89288 15264 89608 16288
rect 89288 15200 89296 15264
rect 89360 15200 89376 15264
rect 89440 15200 89456 15264
rect 89520 15200 89536 15264
rect 89600 15200 89608 15264
rect 89288 14176 89608 15200
rect 89288 14112 89296 14176
rect 89360 14112 89376 14176
rect 89440 14112 89456 14176
rect 89520 14112 89536 14176
rect 89600 14112 89608 14176
rect 89288 13088 89608 14112
rect 89288 13024 89296 13088
rect 89360 13024 89376 13088
rect 89440 13024 89456 13088
rect 89520 13024 89536 13088
rect 89600 13024 89608 13088
rect 89288 12000 89608 13024
rect 89288 11936 89296 12000
rect 89360 11936 89376 12000
rect 89440 11936 89456 12000
rect 89520 11936 89536 12000
rect 89600 11936 89608 12000
rect 89288 10912 89608 11936
rect 89288 10848 89296 10912
rect 89360 10848 89376 10912
rect 89440 10848 89456 10912
rect 89520 10848 89536 10912
rect 89600 10848 89608 10912
rect 89288 9824 89608 10848
rect 89288 9760 89296 9824
rect 89360 9760 89376 9824
rect 89440 9760 89456 9824
rect 89520 9760 89536 9824
rect 89600 9760 89608 9824
rect 89288 8736 89608 9760
rect 89288 8672 89296 8736
rect 89360 8672 89376 8736
rect 89440 8672 89456 8736
rect 89520 8672 89536 8736
rect 89600 8672 89608 8736
rect 89288 7648 89608 8672
rect 89288 7584 89296 7648
rect 89360 7584 89376 7648
rect 89440 7584 89456 7648
rect 89520 7584 89536 7648
rect 89600 7584 89608 7648
rect 89288 6560 89608 7584
rect 89288 6496 89296 6560
rect 89360 6496 89376 6560
rect 89440 6496 89456 6560
rect 89520 6496 89536 6560
rect 89600 6496 89608 6560
rect 89288 5472 89608 6496
rect 89288 5408 89296 5472
rect 89360 5408 89376 5472
rect 89440 5408 89456 5472
rect 89520 5408 89536 5472
rect 89600 5408 89608 5472
rect 89288 4384 89608 5408
rect 89288 4320 89296 4384
rect 89360 4320 89376 4384
rect 89440 4320 89456 4384
rect 89520 4320 89536 4384
rect 89600 4320 89608 4384
rect 89288 3296 89608 4320
rect 89288 3232 89296 3296
rect 89360 3232 89376 3296
rect 89440 3232 89456 3296
rect 89520 3232 89536 3296
rect 89600 3232 89608 3296
rect 89288 2208 89608 3232
rect 89288 2144 89296 2208
rect 89360 2144 89376 2208
rect 89440 2144 89456 2208
rect 89520 2144 89536 2208
rect 89600 2144 89608 2208
rect 89288 2128 89608 2144
rect 104012 27776 104332 27792
rect 104012 27712 104020 27776
rect 104084 27712 104100 27776
rect 104164 27712 104180 27776
rect 104244 27712 104260 27776
rect 104324 27712 104332 27776
rect 104012 26688 104332 27712
rect 104012 26624 104020 26688
rect 104084 26624 104100 26688
rect 104164 26624 104180 26688
rect 104244 26624 104260 26688
rect 104324 26624 104332 26688
rect 104012 25600 104332 26624
rect 104012 25536 104020 25600
rect 104084 25536 104100 25600
rect 104164 25536 104180 25600
rect 104244 25536 104260 25600
rect 104324 25536 104332 25600
rect 104012 24512 104332 25536
rect 104012 24448 104020 24512
rect 104084 24448 104100 24512
rect 104164 24448 104180 24512
rect 104244 24448 104260 24512
rect 104324 24448 104332 24512
rect 104012 23424 104332 24448
rect 104012 23360 104020 23424
rect 104084 23360 104100 23424
rect 104164 23360 104180 23424
rect 104244 23360 104260 23424
rect 104324 23360 104332 23424
rect 104012 22336 104332 23360
rect 104012 22272 104020 22336
rect 104084 22272 104100 22336
rect 104164 22272 104180 22336
rect 104244 22272 104260 22336
rect 104324 22272 104332 22336
rect 104012 21248 104332 22272
rect 104012 21184 104020 21248
rect 104084 21184 104100 21248
rect 104164 21184 104180 21248
rect 104244 21184 104260 21248
rect 104324 21184 104332 21248
rect 104012 20160 104332 21184
rect 104012 20096 104020 20160
rect 104084 20096 104100 20160
rect 104164 20096 104180 20160
rect 104244 20096 104260 20160
rect 104324 20096 104332 20160
rect 104012 19072 104332 20096
rect 104012 19008 104020 19072
rect 104084 19008 104100 19072
rect 104164 19008 104180 19072
rect 104244 19008 104260 19072
rect 104324 19008 104332 19072
rect 104012 17984 104332 19008
rect 104012 17920 104020 17984
rect 104084 17920 104100 17984
rect 104164 17920 104180 17984
rect 104244 17920 104260 17984
rect 104324 17920 104332 17984
rect 104012 16896 104332 17920
rect 104012 16832 104020 16896
rect 104084 16832 104100 16896
rect 104164 16832 104180 16896
rect 104244 16832 104260 16896
rect 104324 16832 104332 16896
rect 104012 15808 104332 16832
rect 104012 15744 104020 15808
rect 104084 15744 104100 15808
rect 104164 15744 104180 15808
rect 104244 15744 104260 15808
rect 104324 15744 104332 15808
rect 104012 14720 104332 15744
rect 104012 14656 104020 14720
rect 104084 14656 104100 14720
rect 104164 14656 104180 14720
rect 104244 14656 104260 14720
rect 104324 14656 104332 14720
rect 104012 13632 104332 14656
rect 104012 13568 104020 13632
rect 104084 13568 104100 13632
rect 104164 13568 104180 13632
rect 104244 13568 104260 13632
rect 104324 13568 104332 13632
rect 104012 12544 104332 13568
rect 104012 12480 104020 12544
rect 104084 12480 104100 12544
rect 104164 12480 104180 12544
rect 104244 12480 104260 12544
rect 104324 12480 104332 12544
rect 104012 11456 104332 12480
rect 104012 11392 104020 11456
rect 104084 11392 104100 11456
rect 104164 11392 104180 11456
rect 104244 11392 104260 11456
rect 104324 11392 104332 11456
rect 104012 10368 104332 11392
rect 104012 10304 104020 10368
rect 104084 10304 104100 10368
rect 104164 10304 104180 10368
rect 104244 10304 104260 10368
rect 104324 10304 104332 10368
rect 104012 9280 104332 10304
rect 104012 9216 104020 9280
rect 104084 9216 104100 9280
rect 104164 9216 104180 9280
rect 104244 9216 104260 9280
rect 104324 9216 104332 9280
rect 104012 8192 104332 9216
rect 104012 8128 104020 8192
rect 104084 8128 104100 8192
rect 104164 8128 104180 8192
rect 104244 8128 104260 8192
rect 104324 8128 104332 8192
rect 104012 7104 104332 8128
rect 104012 7040 104020 7104
rect 104084 7040 104100 7104
rect 104164 7040 104180 7104
rect 104244 7040 104260 7104
rect 104324 7040 104332 7104
rect 104012 6016 104332 7040
rect 104012 5952 104020 6016
rect 104084 5952 104100 6016
rect 104164 5952 104180 6016
rect 104244 5952 104260 6016
rect 104324 5952 104332 6016
rect 104012 4928 104332 5952
rect 104012 4864 104020 4928
rect 104084 4864 104100 4928
rect 104164 4864 104180 4928
rect 104244 4864 104260 4928
rect 104324 4864 104332 4928
rect 104012 3840 104332 4864
rect 104012 3776 104020 3840
rect 104084 3776 104100 3840
rect 104164 3776 104180 3840
rect 104244 3776 104260 3840
rect 104324 3776 104332 3840
rect 104012 2752 104332 3776
rect 104012 2688 104020 2752
rect 104084 2688 104100 2752
rect 104164 2688 104180 2752
rect 104244 2688 104260 2752
rect 104324 2688 104332 2752
rect 104012 2128 104332 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 58696 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1649977179
transform -1 0 85652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1649977179
transform -1 0 33304 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1649977179
transform -1 0 95588 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1649977179
transform 1 0 84088 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1649977179
transform -1 0 76176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1649977179
transform -1 0 59708 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1649977179
transform -1 0 31004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1649977179
transform -1 0 67896 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1649977179
transform 1 0 1840 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1649977179
transform -1 0 117760 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1649977179
transform 1 0 109756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1649977179
transform 1 0 2944 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1649977179
transform -1 0 117760 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1649977179
transform 1 0 1840 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1649977179
transform -1 0 30452 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1649977179
transform -1 0 79856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1649977179
transform 1 0 74244 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1649977179
transform 1 0 28336 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1649977179
transform -1 0 64492 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1649977179
transform -1 0 62744 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1649977179
transform 1 0 12052 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1649977179
transform 1 0 11040 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1649977179
transform 1 0 56304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1649977179
transform 1 0 54832 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1649977179
transform -1 0 107916 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1649977179
transform -1 0 108284 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1649977179
transform -1 0 69000 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1649977179
transform -1 0 38640 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1649977179
transform -1 0 81972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1649977179
transform 1 0 66608 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1649977179
transform 1 0 69184 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1649977179
transform 1 0 67712 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1649977179
transform 1 0 116748 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1649977179
transform 1 0 117668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1649977179
transform 1 0 7452 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1649977179
transform 1 0 71760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1649977179
transform 1 0 68908 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1649977179
transform 1 0 70288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1649977179
transform 1 0 68540 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1649977179
transform 1 0 71208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1649977179
transform 1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1649977179
transform 1 0 76176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1649977179
transform 1 0 30728 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1649977179
transform 1 0 76636 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1649977179
transform 1 0 78016 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1649977179
transform 1 0 24840 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1649977179
transform 1 0 25760 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1649977179
transform 1 0 66516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1649977179
transform 1 0 69736 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1649977179
transform 1 0 79304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1649977179
transform 1 0 72496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1649977179
transform 1 0 90896 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1649977179
transform 1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1649977179
transform 1 0 38088 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_61
timestamp 1649977179
transform 1 0 116840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_62
timestamp 1649977179
transform 1 0 72588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_63
timestamp 1649977179
transform 1 0 53084 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_64
timestamp 1649977179
transform 1 0 100188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_65
timestamp 1649977179
transform 1 0 55476 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_66
timestamp 1649977179
transform 1 0 40848 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_67
timestamp 1649977179
transform 1 0 73508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_68
timestamp 1649977179
transform 1 0 60260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_69
timestamp 1649977179
transform 1 0 41124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_70
timestamp 1649977179
transform 1 0 89700 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_71
timestamp 1649977179
transform 1 0 89332 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_72
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_73
timestamp 1649977179
transform 1 0 36708 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_74
timestamp 1649977179
transform -1 0 83352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_75
timestamp 1649977179
transform 1 0 33120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_76
timestamp 1649977179
transform 1 0 66332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_77
timestamp 1649977179
transform 1 0 31648 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78
timestamp 1649977179
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1649977179
transform 1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95
timestamp 1649977179
transform 1 0 9844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_102
timestamp 1649977179
transform 1 0 10488 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12696 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1649977179
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_172
timestamp 1649977179
transform 1 0 16928 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_200
timestamp 1649977179
transform 1 0 19504 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 1649977179
transform 1 0 19872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1649977179
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1649977179
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 1649977179
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1649977179
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_266
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_272 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_314
timestamp 1649977179
transform 1 0 29992 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_325
timestamp 1649977179
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_346
timestamp 1649977179
transform 1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_350
timestamp 1649977179
transform 1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1649977179
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1649977179
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398
timestamp 1649977179
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_404
timestamp 1649977179
transform 1 0 38272 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_409
timestamp 1649977179
transform 1 0 38732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1649977179
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_421
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_433
timestamp 1649977179
transform 1 0 40940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_437
timestamp 1649977179
transform 1 0 41308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_443
timestamp 1649977179
transform 1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1649977179
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_467
timestamp 1649977179
transform 1 0 44068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1649977179
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_485
timestamp 1649977179
transform 1 0 45724 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_489
timestamp 1649977179
transform 1 0 46092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1649977179
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_514
timestamp 1649977179
transform 1 0 48392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_520
timestamp 1649977179
transform 1 0 48944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_524
timestamp 1649977179
transform 1 0 49312 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_556
timestamp 1649977179
transform 1 0 52256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_570
timestamp 1649977179
transform 1 0 53544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_577
timestamp 1649977179
transform 1 0 54188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_584
timestamp 1649977179
transform 1 0 54832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_589
timestamp 1649977179
transform 1 0 55292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_593
timestamp 1649977179
transform 1 0 55660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_598
timestamp 1649977179
transform 1 0 56120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_612
timestamp 1649977179
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1649977179
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_623
timestamp 1649977179
transform 1 0 58420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_636
timestamp 1649977179
transform 1 0 59616 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_645
timestamp 1649977179
transform 1 0 60444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_656
timestamp 1649977179
transform 1 0 61456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_663
timestamp 1649977179
transform 1 0 62100 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_671
timestamp 1649977179
transform 1 0 62836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_673
timestamp 1649977179
transform 1 0 63020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_678
timestamp 1649977179
transform 1 0 63480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_685
timestamp 1649977179
transform 1 0 64124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_692
timestamp 1649977179
transform 1 0 64768 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_701
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_706
timestamp 1649977179
transform 1 0 66056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_711
timestamp 1649977179
transform 1 0 66516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_722
timestamp 1649977179
transform 1 0 67528 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_735
timestamp 1649977179
transform 1 0 68724 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_739
timestamp 1649977179
transform 1 0 69092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_750
timestamp 1649977179
transform 1 0 70104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_754
timestamp 1649977179
transform 1 0 70472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_760
timestamp 1649977179
transform 1 0 71024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_764
timestamp 1649977179
transform 1 0 71392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_775
timestamp 1649977179
transform 1 0 72404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_779
timestamp 1649977179
transform 1 0 72772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_783
timestamp 1649977179
transform 1 0 73140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_785
timestamp 1649977179
transform 1 0 73324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_793
timestamp 1649977179
transform 1 0 74060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_801
timestamp 1649977179
transform 1 0 74796 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_813
timestamp 1649977179
transform 1 0 75900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_818
timestamp 1649977179
transform 1 0 76360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_829
timestamp 1649977179
transform 1 0 77372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_836
timestamp 1649977179
transform 1 0 78016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_841
timestamp 1649977179
transform 1 0 78476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_846
timestamp 1649977179
transform 1 0 78936 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1649977179
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1649977179
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_879
timestamp 1649977179
transform 1 0 81972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_887
timestamp 1649977179
transform 1 0 82708 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_895
timestamp 1649977179
transform 1 0 83444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_901
timestamp 1649977179
transform 1 0 83996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_908
timestamp 1649977179
transform 1 0 84640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_912
timestamp 1649977179
transform 1 0 85008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_916
timestamp 1649977179
transform 1 0 85376 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_928
timestamp 1649977179
transform 1 0 86480 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_936
timestamp 1649977179
transform 1 0 87216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_948
timestamp 1649977179
transform 1 0 88320 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_956
timestamp 1649977179
transform 1 0 89056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_965
timestamp 1649977179
transform 1 0 89884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_972
timestamp 1649977179
transform 1 0 90528 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_981
timestamp 1649977179
transform 1 0 91356 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_986
timestamp 1649977179
transform 1 0 91816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_993
timestamp 1649977179
transform 1 0 92460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1001
timestamp 1649977179
transform 1 0 93196 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1007
timestamp 1649977179
transform 1 0 93748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1009
timestamp 1649977179
transform 1 0 93932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1014
timestamp 1649977179
transform 1 0 94392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1024
timestamp 1649977179
transform 1 0 95312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1028
timestamp 1649977179
transform 1 0 95680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1032
timestamp 1649977179
transform 1 0 96048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1037
timestamp 1649977179
transform 1 0 96508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1045
timestamp 1649977179
transform 1 0 97244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1057
timestamp 1649977179
transform 1 0 98348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1063
timestamp 1649977179
transform 1 0 98900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1065
timestamp 1649977179
transform 1 0 99084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1073
timestamp 1649977179
transform 1 0 99820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1079
timestamp 1649977179
transform 1 0 100372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1085
timestamp 1649977179
transform 1 0 100924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1091
timestamp 1649977179
transform 1 0 101476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1093
timestamp 1649977179
transform 1 0 101660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1103
timestamp 1649977179
transform 1 0 102580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1113
timestamp 1649977179
transform 1 0 103500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1119
timestamp 1649977179
transform 1 0 104052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1121
timestamp 1649977179
transform 1 0 104236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1126
timestamp 1649977179
transform 1 0 104696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1134
timestamp 1649977179
transform 1 0 105432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1141
timestamp 1649977179
transform 1 0 106076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1147
timestamp 1649977179
transform 1 0 106628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1152
timestamp 1649977179
transform 1 0 107088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1159
timestamp 1649977179
transform 1 0 107732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1166
timestamp 1649977179
transform 1 0 108376 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1174
timestamp 1649977179
transform 1 0 109112 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1177
timestamp 1649977179
transform 1 0 109388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1185
timestamp 1649977179
transform 1 0 110124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1197
timestamp 1649977179
transform 1 0 111228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1203
timestamp 1649977179
transform 1 0 111780 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1205
timestamp 1649977179
transform 1 0 111964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1217
timestamp 1649977179
transform 1 0 113068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1224
timestamp 1649977179
transform 1 0 113712 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1236
timestamp 1649977179
transform 1 0 114816 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1246
timestamp 1649977179
transform 1 0 115736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1256
timestamp 1649977179
transform 1 0 116656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1261
timestamp 1649977179
transform 1 0 117116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1271
timestamp 1649977179
transform 1 0 118036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_18
timestamp 1649977179
transform 1 0 2760 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_22
timestamp 1649977179
transform 1 0 3128 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1649977179
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_60
timestamp 1649977179
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_64
timestamp 1649977179
transform 1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_80
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_92
timestamp 1649977179
transform 1 0 9568 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_102
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_122
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_134
timestamp 1649977179
transform 1 0 13432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1649977179
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_146
timestamp 1649977179
transform 1 0 14536 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1649977179
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1649977179
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_267
timestamp 1649977179
transform 1 0 25668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1649977179
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1649977179
transform 1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_304
timestamp 1649977179
transform 1 0 29072 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_312
timestamp 1649977179
transform 1 0 29808 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_324
timestamp 1649977179
transform 1 0 30912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_328
timestamp 1649977179
transform 1 0 31280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_347
timestamp 1649977179
transform 1 0 33028 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_354
timestamp 1649977179
transform 1 0 33672 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_366
timestamp 1649977179
transform 1 0 34776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1649977179
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_378
timestamp 1649977179
transform 1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_413
timestamp 1649977179
transform 1 0 39100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1649977179
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_432
timestamp 1649977179
transform 1 0 40848 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_440
timestamp 1649977179
transform 1 0 41584 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1649977179
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_460
timestamp 1649977179
transform 1 0 43424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_464
timestamp 1649977179
transform 1 0 43792 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_468
timestamp 1649977179
transform 1 0 44160 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_484
timestamp 1649977179
transform 1 0 45632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_492
timestamp 1649977179
transform 1 0 46368 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1649977179
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_510
timestamp 1649977179
transform 1 0 48024 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1649977179
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_541
timestamp 1649977179
transform 1 0 50876 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_545
timestamp 1649977179
transform 1 0 51244 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_555
timestamp 1649977179
transform 1 0 52164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1649977179
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1649977179
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_566
timestamp 1649977179
transform 1 0 53176 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_578
timestamp 1649977179
transform 1 0 54280 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_590
timestamp 1649977179
transform 1 0 55384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_594
timestamp 1649977179
transform 1 0 55752 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_602
timestamp 1649977179
transform 1 0 56488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_612
timestamp 1649977179
transform 1 0 57408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_621
timestamp 1649977179
transform 1 0 58236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_630
timestamp 1649977179
transform 1 0 59064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_644
timestamp 1649977179
transform 1 0 60352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_652
timestamp 1649977179
transform 1 0 61088 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_660
timestamp 1649977179
transform 1 0 61824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_664
timestamp 1649977179
transform 1 0 62192 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1649977179
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_685
timestamp 1649977179
transform 1 0 64124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_691
timestamp 1649977179
transform 1 0 64676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_698
timestamp 1649977179
transform 1 0 65320 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_706
timestamp 1649977179
transform 1 0 66056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_710
timestamp 1649977179
transform 1 0 66424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_717
timestamp 1649977179
transform 1 0 67068 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_725
timestamp 1649977179
transform 1 0 67804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_729
timestamp 1649977179
transform 1 0 68172 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_734
timestamp 1649977179
transform 1 0 68632 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_742
timestamp 1649977179
transform 1 0 69368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_748
timestamp 1649977179
transform 1 0 69920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_756
timestamp 1649977179
transform 1 0 70656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_760
timestamp 1649977179
transform 1 0 71024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_765
timestamp 1649977179
transform 1 0 71484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_778
timestamp 1649977179
transform 1 0 72680 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_788
timestamp 1649977179
transform 1 0 73600 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_796
timestamp 1649977179
transform 1 0 74336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_801
timestamp 1649977179
transform 1 0 74796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_809
timestamp 1649977179
transform 1 0 75532 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_817
timestamp 1649977179
transform 1 0 76268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_828
timestamp 1649977179
transform 1 0 77280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_835
timestamp 1649977179
transform 1 0 77924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1649977179
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1649977179
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1649977179
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_865
timestamp 1649977179
transform 1 0 80684 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_874
timestamp 1649977179
transform 1 0 81512 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_886
timestamp 1649977179
transform 1 0 82616 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_894
timestamp 1649977179
transform 1 0 83352 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1649977179
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1649977179
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1649977179
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_933
timestamp 1649977179
transform 1 0 86940 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_937
timestamp 1649977179
transform 1 0 87308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_949
timestamp 1649977179
transform 1 0 88412 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1649977179
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1649977179
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1649977179
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1649977179
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1649977179
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1649977179
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1649977179
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1649977179
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1649977179
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1649977179
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1649977179
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1649977179
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1068
timestamp 1649977179
transform 1 0 99360 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1080
timestamp 1649977179
transform 1 0 100464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1092
timestamp 1649977179
transform 1 0 101568 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1100
timestamp 1649977179
transform 1 0 102304 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1105
timestamp 1649977179
transform 1 0 102764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1117
timestamp 1649977179
transform 1 0 103868 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1649977179
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1649977179
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1145
timestamp 1649977179
transform 1 0 106444 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1153
timestamp 1649977179
transform 1 0 107180 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1159
timestamp 1649977179
transform 1 0 107732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1171
timestamp 1649977179
transform 1 0 108836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1649977179
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1177
timestamp 1649977179
transform 1 0 109388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1183
timestamp 1649977179
transform 1 0 109940 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1188
timestamp 1649977179
transform 1 0 110400 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1204
timestamp 1649977179
transform 1 0 111872 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1216
timestamp 1649977179
transform 1 0 112976 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1228
timestamp 1649977179
transform 1 0 114080 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1233
timestamp 1649977179
transform 1 0 114540 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1245
timestamp 1649977179
transform 1 0 115644 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1252
timestamp 1649977179
transform 1 0 116288 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1258
timestamp 1649977179
transform 1 0 116840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1263
timestamp 1649977179
transform 1 0 117300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1273
timestamp 1649977179
transform 1 0 118220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_6
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1649977179
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_341
timestamp 1649977179
transform 1 0 32476 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_346
timestamp 1649977179
transform 1 0 32936 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_358
timestamp 1649977179
transform 1 0 34040 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_429
timestamp 1649977179
transform 1 0 40572 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_454
timestamp 1649977179
transform 1 0 42872 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_466
timestamp 1649977179
transform 1 0 43976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1649977179
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_485
timestamp 1649977179
transform 1 0 45724 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_500
timestamp 1649977179
transform 1 0 47104 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_507
timestamp 1649977179
transform 1 0 47748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_519
timestamp 1649977179
transform 1 0 48852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_553
timestamp 1649977179
transform 1 0 51980 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_559
timestamp 1649977179
transform 1 0 52532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_571
timestamp 1649977179
transform 1 0 53636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_583
timestamp 1649977179
transform 1 0 54740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1649977179
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_601
timestamp 1649977179
transform 1 0 56396 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_609
timestamp 1649977179
transform 1 0 57132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_615
timestamp 1649977179
transform 1 0 57684 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_622
timestamp 1649977179
transform 1 0 58328 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_638
timestamp 1649977179
transform 1 0 59800 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_645
timestamp 1649977179
transform 1 0 60444 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_653
timestamp 1649977179
transform 1 0 61180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_665
timestamp 1649977179
transform 1 0 62284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_677
timestamp 1649977179
transform 1 0 63388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_689
timestamp 1649977179
transform 1 0 64492 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_697
timestamp 1649977179
transform 1 0 65228 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1649977179
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1649977179
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1649977179
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1649977179
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_760
timestamp 1649977179
transform 1 0 71024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_767
timestamp 1649977179
transform 1 0 71668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_774
timestamp 1649977179
transform 1 0 72312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_778
timestamp 1649977179
transform 1 0 72680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_783
timestamp 1649977179
transform 1 0 73140 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_791
timestamp 1649977179
transform 1 0 73876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_795
timestamp 1649977179
transform 1 0 74244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_804
timestamp 1649977179
transform 1 0 75072 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_816
timestamp 1649977179
transform 1 0 76176 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_828
timestamp 1649977179
transform 1 0 77280 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_840
timestamp 1649977179
transform 1 0 78384 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_852
timestamp 1649977179
transform 1 0 79488 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_864
timestamp 1649977179
transform 1 0 80592 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1649977179
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1649977179
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1649977179
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1649977179
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1649977179
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1649977179
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1649977179
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1649977179
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1649977179
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1649977179
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1649977179
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1649977179
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1649977179
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1649977179
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1649977179
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1649977179
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1649977179
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1649977179
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1649977179
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1649977179
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1649977179
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1649977179
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1649977179
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1649977179
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1649977179
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1649977179
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1649977179
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1649977179
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1649977179
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1649977179
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1649977179
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1649977179
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1649977179
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1185
timestamp 1649977179
transform 1 0 110124 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1197
timestamp 1649977179
transform 1 0 111228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1649977179
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1649977179
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1217
timestamp 1649977179
transform 1 0 113068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1229
timestamp 1649977179
transform 1 0 114172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1241
timestamp 1649977179
transform 1 0 115276 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1256
timestamp 1649977179
transform 1 0 116656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1261
timestamp 1649977179
transform 1 0 117116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1265
timestamp 1649977179
transform 1 0 117484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1273
timestamp 1649977179
transform 1 0 118220 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6
timestamp 1649977179
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_18
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_30
timestamp 1649977179
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_42
timestamp 1649977179
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_629
timestamp 1649977179
transform 1 0 58972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_636
timestamp 1649977179
transform 1 0 59616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_642
timestamp 1649977179
transform 1 0 60168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_645
timestamp 1649977179
transform 1 0 60444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_656
timestamp 1649977179
transform 1 0 61456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_663
timestamp 1649977179
transform 1 0 62100 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1649977179
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1649977179
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1649977179
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1649977179
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1649977179
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1649977179
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1649977179
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1649977179
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1649977179
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1649977179
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1649977179
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1649977179
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1649977179
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1649977179
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_841
timestamp 1649977179
transform 1 0 78476 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_850
timestamp 1649977179
transform 1 0 79304 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_862
timestamp 1649977179
transform 1 0 80408 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_874
timestamp 1649977179
transform 1 0 81512 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_880
timestamp 1649977179
transform 1 0 82064 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_890
timestamp 1649977179
transform 1 0 82984 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1649977179
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1649977179
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1649977179
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1649977179
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1649977179
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1649977179
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1649977179
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1649977179
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1649977179
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1649977179
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1649977179
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1649977179
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1649977179
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1649977179
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1649977179
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1649977179
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1649977179
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1649977179
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1649977179
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1649977179
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1649977179
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1649977179
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1649977179
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1649977179
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1649977179
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1649977179
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1649977179
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1649977179
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1649977179
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1649977179
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1649977179
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1649977179
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1649977179
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1649977179
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1649977179
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1649977179
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1649977179
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1649977179
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1257
timestamp 1649977179
transform 1 0 116748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1260
timestamp 1649977179
transform 1 0 117024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1265
timestamp 1649977179
transform 1 0 117484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1273
timestamp 1649977179
transform 1 0 118220 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1649977179
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1649977179
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1649977179
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1649977179
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1649977179
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1649977179
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1649977179
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1649977179
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1649977179
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1649977179
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1649977179
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1649977179
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1649977179
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1649977179
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1649977179
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1649977179
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1649977179
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1649977179
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1649977179
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1649977179
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1649977179
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1649977179
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1649977179
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_849
timestamp 1649977179
transform 1 0 79212 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_852
timestamp 1649977179
transform 1 0 79488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_858
timestamp 1649977179
transform 1 0 80040 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_866
timestamp 1649977179
transform 1 0 80776 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1649977179
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1649977179
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1649977179
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1649977179
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1649977179
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1649977179
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1649977179
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1649977179
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1649977179
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1649977179
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1649977179
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1649977179
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1649977179
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1649977179
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1649977179
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1649977179
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1649977179
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1649977179
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1649977179
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1649977179
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1649977179
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1649977179
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1649977179
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1649977179
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1649977179
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1649977179
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1649977179
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1649977179
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1649977179
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1649977179
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1649977179
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1649977179
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1649977179
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1649977179
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1649977179
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1649977179
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1649977179
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1217
timestamp 1649977179
transform 1 0 113068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1229
timestamp 1649977179
transform 1 0 114172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1241
timestamp 1649977179
transform 1 0 115276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1253
timestamp 1649977179
transform 1 0 116380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1649977179
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1261
timestamp 1649977179
transform 1 0 117116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1273
timestamp 1649977179
transform 1 0 118220 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1649977179
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1649977179
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1649977179
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1649977179
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1649977179
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1649977179
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1649977179
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1649977179
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1649977179
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1649977179
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1649977179
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1649977179
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1649977179
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1649977179
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1649977179
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1649977179
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1649977179
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1649977179
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1649977179
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1649977179
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_877
timestamp 1649977179
transform 1 0 81788 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_885
timestamp 1649977179
transform 1 0 82524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_891
timestamp 1649977179
transform 1 0 83076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1649977179
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1649977179
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1649977179
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1649977179
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1649977179
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1649977179
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1649977179
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1649977179
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1649977179
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1649977179
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1649977179
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1649977179
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1649977179
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1649977179
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1649977179
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1649977179
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1649977179
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1649977179
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1649977179
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1649977179
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1649977179
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1649977179
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1649977179
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1649977179
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1649977179
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1649977179
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1649977179
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1649977179
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1649977179
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1649977179
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1649977179
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1649977179
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1649977179
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1649977179
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1649977179
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1649977179
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1649977179
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1649977179
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1245
timestamp 1649977179
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1257
timestamp 1649977179
transform 1 0 116748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1269
timestamp 1649977179
transform 1 0 117852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1273
timestamp 1649977179
transform 1 0 118220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_11
timestamp 1649977179
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1649977179
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1649977179
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1649977179
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1649977179
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1649977179
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1649977179
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1649977179
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1649977179
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1649977179
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1649977179
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1649977179
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1649977179
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1649977179
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1649977179
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1649977179
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1649977179
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1649977179
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1649977179
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1649977179
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1649977179
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1649977179
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1649977179
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1649977179
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1649977179
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1649977179
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1649977179
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1649977179
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1649977179
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1649977179
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1649977179
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1649977179
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1649977179
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1649977179
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1649977179
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1649977179
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1649977179
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1649977179
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1649977179
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1649977179
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1649977179
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1649977179
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1649977179
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1649977179
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1649977179
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1649977179
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1649977179
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1649977179
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1649977179
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1649977179
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1649977179
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1649977179
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1649977179
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1649977179
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1649977179
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1649977179
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1649977179
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1649977179
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1229
timestamp 1649977179
transform 1 0 114172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1241
timestamp 1649977179
transform 1 0 115276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1649977179
transform 1 0 116380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1649977179
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1261
timestamp 1649977179
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1273
timestamp 1649977179
transform 1 0 118220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_10
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_22
timestamp 1649977179
transform 1 0 3128 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_34
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1649977179
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_539
timestamp 1649977179
transform 1 0 50692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_551
timestamp 1649977179
transform 1 0 51796 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1649977179
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1649977179
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1649977179
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1649977179
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1649977179
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1649977179
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1649977179
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1649977179
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1649977179
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1649977179
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1649977179
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1649977179
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1649977179
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1649977179
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1649977179
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1649977179
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1649977179
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1649977179
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1649977179
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1649977179
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_921
timestamp 1649977179
transform 1 0 85836 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_929
timestamp 1649977179
transform 1 0 86572 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_934
timestamp 1649977179
transform 1 0 87032 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_946
timestamp 1649977179
transform 1 0 88136 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1649977179
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1649977179
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1649977179
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1649977179
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1649977179
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1649977179
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1649977179
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1649977179
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1649977179
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1649977179
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1649977179
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1649977179
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1649977179
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1649977179
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1649977179
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1649977179
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1649977179
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1649977179
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1649977179
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1649977179
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1649977179
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1649977179
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1649977179
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1649977179
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1649977179
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1189
timestamp 1649977179
transform 1 0 110492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1201
timestamp 1649977179
transform 1 0 111596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1213
timestamp 1649977179
transform 1 0 112700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1649977179
transform 1 0 113804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1649977179
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1233
timestamp 1649977179
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1245
timestamp 1649977179
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1257
timestamp 1649977179
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1273
timestamp 1649977179
transform 1 0 118220 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_536
timestamp 1649977179
transform 1 0 50416 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_548
timestamp 1649977179
transform 1 0 51520 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_560
timestamp 1649977179
transform 1 0 52624 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_572
timestamp 1649977179
transform 1 0 53728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_584
timestamp 1649977179
transform 1 0 54832 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1649977179
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1649977179
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1649977179
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1649977179
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1649977179
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1649977179
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1649977179
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1649977179
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1649977179
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1649977179
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1649977179
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1649977179
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1649977179
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1649977179
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1649977179
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1649977179
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1649977179
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1649977179
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1649977179
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1649977179
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1649977179
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1649977179
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1649977179
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1649977179
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1649977179
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1649977179
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1649977179
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1649977179
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1649977179
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1649977179
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1649977179
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1649977179
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1649977179
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1649977179
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1649977179
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1649977179
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1649977179
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1649977179
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1649977179
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1649977179
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1649977179
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1649977179
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1649977179
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1649977179
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1649977179
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1649977179
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1649977179
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1649977179
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1649977179
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1161
timestamp 1649977179
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1649977179
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1185
timestamp 1649977179
transform 1 0 110124 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1649977179
transform 1 0 111228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1649977179
transform 1 0 111780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1205
timestamp 1649977179
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1217
timestamp 1649977179
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1229
timestamp 1649977179
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1241
timestamp 1649977179
transform 1 0 115276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1649977179
transform 1 0 116380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1649977179
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1261
timestamp 1649977179
transform 1 0 117116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1273
timestamp 1649977179
transform 1 0 118220 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1649977179
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1649977179
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1649977179
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1649977179
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1649977179
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1649977179
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1649977179
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1649977179
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_821
timestamp 1649977179
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1649977179
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1649977179
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1649977179
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1649977179
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_865
timestamp 1649977179
transform 1 0 80684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_877
timestamp 1649977179
transform 1 0 81788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_889
timestamp 1649977179
transform 1 0 82892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_895
timestamp 1649977179
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1649977179
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1649977179
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_921
timestamp 1649977179
transform 1 0 85836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_930
timestamp 1649977179
transform 1 0 86664 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_942
timestamp 1649977179
transform 1 0 87768 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_950
timestamp 1649977179
transform 1 0 88504 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1649977179
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1649977179
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_977
timestamp 1649977179
transform 1 0 90988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_989
timestamp 1649977179
transform 1 0 92092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1001
timestamp 1649977179
transform 1 0 93196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1007
timestamp 1649977179
transform 1 0 93748 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1649977179
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1649977179
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1033
timestamp 1649977179
transform 1 0 96140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1045
timestamp 1649977179
transform 1 0 97244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1057
timestamp 1649977179
transform 1 0 98348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1063
timestamp 1649977179
transform 1 0 98900 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1649977179
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1649977179
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1089
timestamp 1649977179
transform 1 0 101292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1101
timestamp 1649977179
transform 1 0 102396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1113
timestamp 1649977179
transform 1 0 103500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1119
timestamp 1649977179
transform 1 0 104052 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1649977179
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1649977179
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1145
timestamp 1649977179
transform 1 0 106444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1157
timestamp 1649977179
transform 1 0 107548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1169
timestamp 1649977179
transform 1 0 108652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1175
timestamp 1649977179
transform 1 0 109204 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1649977179
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1189
timestamp 1649977179
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1201
timestamp 1649977179
transform 1 0 111596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1213
timestamp 1649977179
transform 1 0 112700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1225
timestamp 1649977179
transform 1 0 113804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1231
timestamp 1649977179
transform 1 0 114356 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1649977179
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1649977179
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1257
timestamp 1649977179
transform 1 0 116748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1273
timestamp 1649977179
transform 1 0 118220 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 1649977179
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1649977179
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_320
timestamp 1649977179
transform 1 0 30544 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_324
timestamp 1649977179
transform 1 0 30912 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_336
timestamp 1649977179
transform 1 0 32016 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_348
timestamp 1649977179
transform 1 0 33120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1649977179
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1649977179
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1649977179
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1649977179
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1649977179
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1649977179
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1649977179
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1649977179
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1649977179
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1649977179
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_813
timestamp 1649977179
transform 1 0 75900 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_821
timestamp 1649977179
transform 1 0 76636 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_828
timestamp 1649977179
transform 1 0 77280 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_840
timestamp 1649977179
transform 1 0 78384 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_852
timestamp 1649977179
transform 1 0 79488 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_864
timestamp 1649977179
transform 1 0 80592 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_869
timestamp 1649977179
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_881
timestamp 1649977179
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_893
timestamp 1649977179
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_905
timestamp 1649977179
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_917
timestamp 1649977179
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_923
timestamp 1649977179
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_925
timestamp 1649977179
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_937
timestamp 1649977179
transform 1 0 87308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_949
timestamp 1649977179
transform 1 0 88412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_961
timestamp 1649977179
transform 1 0 89516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_973
timestamp 1649977179
transform 1 0 90620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_979
timestamp 1649977179
transform 1 0 91172 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_981
timestamp 1649977179
transform 1 0 91356 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_993
timestamp 1649977179
transform 1 0 92460 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1005
timestamp 1649977179
transform 1 0 93564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1017
timestamp 1649977179
transform 1 0 94668 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1029
timestamp 1649977179
transform 1 0 95772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1035
timestamp 1649977179
transform 1 0 96324 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1037
timestamp 1649977179
transform 1 0 96508 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1049
timestamp 1649977179
transform 1 0 97612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1061
timestamp 1649977179
transform 1 0 98716 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1073
timestamp 1649977179
transform 1 0 99820 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1085
timestamp 1649977179
transform 1 0 100924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1091
timestamp 1649977179
transform 1 0 101476 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1093
timestamp 1649977179
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1105
timestamp 1649977179
transform 1 0 102764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1117
timestamp 1649977179
transform 1 0 103868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1129
timestamp 1649977179
transform 1 0 104972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1141
timestamp 1649977179
transform 1 0 106076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1147
timestamp 1649977179
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1149
timestamp 1649977179
transform 1 0 106812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1161
timestamp 1649977179
transform 1 0 107916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1173
timestamp 1649977179
transform 1 0 109020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1185
timestamp 1649977179
transform 1 0 110124 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1197
timestamp 1649977179
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1203
timestamp 1649977179
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1205
timestamp 1649977179
transform 1 0 111964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1217
timestamp 1649977179
transform 1 0 113068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1229
timestamp 1649977179
transform 1 0 114172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1241
timestamp 1649977179
transform 1 0 115276 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1253
timestamp 1649977179
transform 1 0 116380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1259
timestamp 1649977179
transform 1 0 116932 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1261
timestamp 1649977179
transform 1 0 117116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1273
timestamp 1649977179
transform 1 0 118220 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_6
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_18
timestamp 1649977179
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_30
timestamp 1649977179
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_42
timestamp 1649977179
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_318
timestamp 1649977179
transform 1 0 30360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1649977179
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1649977179
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1649977179
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1649977179
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1649977179
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1649977179
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1649977179
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1649977179
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1649977179
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1649977179
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_821
timestamp 1649977179
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1649977179
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1649977179
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_841
timestamp 1649977179
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_853
timestamp 1649977179
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_865
timestamp 1649977179
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_877
timestamp 1649977179
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1649977179
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1649977179
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_897
timestamp 1649977179
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_909
timestamp 1649977179
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_921
timestamp 1649977179
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_933
timestamp 1649977179
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_945
timestamp 1649977179
transform 1 0 88044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1649977179
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_953
timestamp 1649977179
transform 1 0 88780 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_965
timestamp 1649977179
transform 1 0 89884 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_977
timestamp 1649977179
transform 1 0 90988 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_989
timestamp 1649977179
transform 1 0 92092 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1001
timestamp 1649977179
transform 1 0 93196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1007
timestamp 1649977179
transform 1 0 93748 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1009
timestamp 1649977179
transform 1 0 93932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1021
timestamp 1649977179
transform 1 0 95036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1033
timestamp 1649977179
transform 1 0 96140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1045
timestamp 1649977179
transform 1 0 97244 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1057
timestamp 1649977179
transform 1 0 98348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1063
timestamp 1649977179
transform 1 0 98900 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1065
timestamp 1649977179
transform 1 0 99084 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1077
timestamp 1649977179
transform 1 0 100188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1089
timestamp 1649977179
transform 1 0 101292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1101
timestamp 1649977179
transform 1 0 102396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1113
timestamp 1649977179
transform 1 0 103500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1119
timestamp 1649977179
transform 1 0 104052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1121
timestamp 1649977179
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1133
timestamp 1649977179
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1145
timestamp 1649977179
transform 1 0 106444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1157
timestamp 1649977179
transform 1 0 107548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1169
timestamp 1649977179
transform 1 0 108652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1175
timestamp 1649977179
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1177
timestamp 1649977179
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1189
timestamp 1649977179
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1201
timestamp 1649977179
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1213
timestamp 1649977179
transform 1 0 112700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1225
timestamp 1649977179
transform 1 0 113804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1231
timestamp 1649977179
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1233
timestamp 1649977179
transform 1 0 114540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1245
timestamp 1649977179
transform 1 0 115644 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1257
timestamp 1649977179
transform 1 0 116748 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1265
timestamp 1649977179
transform 1 0 117484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1268
timestamp 1649977179
transform 1 0 117760 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1273
timestamp 1649977179
transform 1 0 118220 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1649977179
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1649977179
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1649977179
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1649977179
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1649977179
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1649977179
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1649977179
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1649977179
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1649977179
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1649977179
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1649977179
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1649977179
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_813
timestamp 1649977179
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_825
timestamp 1649977179
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_837
timestamp 1649977179
transform 1 0 78108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_849
timestamp 1649977179
transform 1 0 79212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_861
timestamp 1649977179
transform 1 0 80316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_867
timestamp 1649977179
transform 1 0 80868 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_869
timestamp 1649977179
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_881
timestamp 1649977179
transform 1 0 82156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_893
timestamp 1649977179
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_905
timestamp 1649977179
transform 1 0 84364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1649977179
transform 1 0 85468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1649977179
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_925
timestamp 1649977179
transform 1 0 86204 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_937
timestamp 1649977179
transform 1 0 87308 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_949
timestamp 1649977179
transform 1 0 88412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_961
timestamp 1649977179
transform 1 0 89516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_973
timestamp 1649977179
transform 1 0 90620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_979
timestamp 1649977179
transform 1 0 91172 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_981
timestamp 1649977179
transform 1 0 91356 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_993
timestamp 1649977179
transform 1 0 92460 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1005
timestamp 1649977179
transform 1 0 93564 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1017
timestamp 1649977179
transform 1 0 94668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1029
timestamp 1649977179
transform 1 0 95772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1035
timestamp 1649977179
transform 1 0 96324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1037
timestamp 1649977179
transform 1 0 96508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1049
timestamp 1649977179
transform 1 0 97612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1061
timestamp 1649977179
transform 1 0 98716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1073
timestamp 1649977179
transform 1 0 99820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1085
timestamp 1649977179
transform 1 0 100924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1091
timestamp 1649977179
transform 1 0 101476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1093
timestamp 1649977179
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1105
timestamp 1649977179
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1117
timestamp 1649977179
transform 1 0 103868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1129
timestamp 1649977179
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1141
timestamp 1649977179
transform 1 0 106076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1147
timestamp 1649977179
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1149
timestamp 1649977179
transform 1 0 106812 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1161
timestamp 1649977179
transform 1 0 107916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1173
timestamp 1649977179
transform 1 0 109020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1185
timestamp 1649977179
transform 1 0 110124 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1197
timestamp 1649977179
transform 1 0 111228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1203
timestamp 1649977179
transform 1 0 111780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1205
timestamp 1649977179
transform 1 0 111964 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1217
timestamp 1649977179
transform 1 0 113068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1229
timestamp 1649977179
transform 1 0 114172 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1241
timestamp 1649977179
transform 1 0 115276 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1253
timestamp 1649977179
transform 1 0 116380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1259
timestamp 1649977179
transform 1 0 116932 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1261
timestamp 1649977179
transform 1 0 117116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1273
timestamp 1649977179
transform 1 0 118220 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1649977179
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1649977179
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1649977179
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1649977179
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1649977179
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1649977179
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1649977179
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1649977179
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1649977179
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1649977179
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1649977179
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1649977179
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1649977179
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1649977179
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1649977179
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_821
timestamp 1649977179
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1649977179
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1649977179
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_841
timestamp 1649977179
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_853
timestamp 1649977179
transform 1 0 79580 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_865
timestamp 1649977179
transform 1 0 80684 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_877
timestamp 1649977179
transform 1 0 81788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_889
timestamp 1649977179
transform 1 0 82892 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_895
timestamp 1649977179
transform 1 0 83444 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_897
timestamp 1649977179
transform 1 0 83628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_909
timestamp 1649977179
transform 1 0 84732 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_921
timestamp 1649977179
transform 1 0 85836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_933
timestamp 1649977179
transform 1 0 86940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_945
timestamp 1649977179
transform 1 0 88044 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_951
timestamp 1649977179
transform 1 0 88596 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_953
timestamp 1649977179
transform 1 0 88780 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_965
timestamp 1649977179
transform 1 0 89884 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_977
timestamp 1649977179
transform 1 0 90988 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_989
timestamp 1649977179
transform 1 0 92092 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1001
timestamp 1649977179
transform 1 0 93196 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1007
timestamp 1649977179
transform 1 0 93748 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1009
timestamp 1649977179
transform 1 0 93932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1021
timestamp 1649977179
transform 1 0 95036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1033
timestamp 1649977179
transform 1 0 96140 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1045
timestamp 1649977179
transform 1 0 97244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1057
timestamp 1649977179
transform 1 0 98348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1063
timestamp 1649977179
transform 1 0 98900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1065
timestamp 1649977179
transform 1 0 99084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1077
timestamp 1649977179
transform 1 0 100188 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1089
timestamp 1649977179
transform 1 0 101292 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1101
timestamp 1649977179
transform 1 0 102396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1113
timestamp 1649977179
transform 1 0 103500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1119
timestamp 1649977179
transform 1 0 104052 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1121
timestamp 1649977179
transform 1 0 104236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1133
timestamp 1649977179
transform 1 0 105340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1145
timestamp 1649977179
transform 1 0 106444 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1157
timestamp 1649977179
transform 1 0 107548 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1169
timestamp 1649977179
transform 1 0 108652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1175
timestamp 1649977179
transform 1 0 109204 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1177
timestamp 1649977179
transform 1 0 109388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1189
timestamp 1649977179
transform 1 0 110492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1201
timestamp 1649977179
transform 1 0 111596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1213
timestamp 1649977179
transform 1 0 112700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1225
timestamp 1649977179
transform 1 0 113804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1231
timestamp 1649977179
transform 1 0 114356 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1236
timestamp 1649977179
transform 1 0 114816 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1248
timestamp 1649977179
transform 1 0 115920 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1260
timestamp 1649977179
transform 1 0 117024 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1272
timestamp 1649977179
transform 1 0 118128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1276
timestamp 1649977179
transform 1 0 118496 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_18
timestamp 1649977179
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1649977179
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1649977179
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1649977179
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1649977179
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1649977179
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1649977179
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1649977179
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1649977179
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1649977179
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1649977179
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1649977179
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1649977179
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1649977179
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1649977179
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1649977179
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_813
timestamp 1649977179
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_825
timestamp 1649977179
transform 1 0 77004 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_837
timestamp 1649977179
transform 1 0 78108 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_849
timestamp 1649977179
transform 1 0 79212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_861
timestamp 1649977179
transform 1 0 80316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_867
timestamp 1649977179
transform 1 0 80868 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_869
timestamp 1649977179
transform 1 0 81052 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_881
timestamp 1649977179
transform 1 0 82156 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_893
timestamp 1649977179
transform 1 0 83260 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_905
timestamp 1649977179
transform 1 0 84364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_917
timestamp 1649977179
transform 1 0 85468 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_923
timestamp 1649977179
transform 1 0 86020 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_925
timestamp 1649977179
transform 1 0 86204 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_937
timestamp 1649977179
transform 1 0 87308 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_949
timestamp 1649977179
transform 1 0 88412 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_961
timestamp 1649977179
transform 1 0 89516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_973
timestamp 1649977179
transform 1 0 90620 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_979
timestamp 1649977179
transform 1 0 91172 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_981
timestamp 1649977179
transform 1 0 91356 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_993
timestamp 1649977179
transform 1 0 92460 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1005
timestamp 1649977179
transform 1 0 93564 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1017
timestamp 1649977179
transform 1 0 94668 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1029
timestamp 1649977179
transform 1 0 95772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1035
timestamp 1649977179
transform 1 0 96324 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1037
timestamp 1649977179
transform 1 0 96508 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1049
timestamp 1649977179
transform 1 0 97612 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1061
timestamp 1649977179
transform 1 0 98716 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1073
timestamp 1649977179
transform 1 0 99820 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1085
timestamp 1649977179
transform 1 0 100924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1091
timestamp 1649977179
transform 1 0 101476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1093
timestamp 1649977179
transform 1 0 101660 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1105
timestamp 1649977179
transform 1 0 102764 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1117
timestamp 1649977179
transform 1 0 103868 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1129
timestamp 1649977179
transform 1 0 104972 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1141
timestamp 1649977179
transform 1 0 106076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1147
timestamp 1649977179
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1149
timestamp 1649977179
transform 1 0 106812 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1161
timestamp 1649977179
transform 1 0 107916 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1173
timestamp 1649977179
transform 1 0 109020 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1185
timestamp 1649977179
transform 1 0 110124 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1197
timestamp 1649977179
transform 1 0 111228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1203
timestamp 1649977179
transform 1 0 111780 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1205
timestamp 1649977179
transform 1 0 111964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1217
timestamp 1649977179
transform 1 0 113068 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1221
timestamp 1649977179
transform 1 0 113436 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1226
timestamp 1649977179
transform 1 0 113896 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1238
timestamp 1649977179
transform 1 0 115000 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1250
timestamp 1649977179
transform 1 0 116104 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1258
timestamp 1649977179
transform 1 0 116840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1261
timestamp 1649977179
transform 1 0 117116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1269
timestamp 1649977179
transform 1 0 117852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1273
timestamp 1649977179
transform 1 0 118220 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_6
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_18
timestamp 1649977179
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_30
timestamp 1649977179
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_42
timestamp 1649977179
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1649977179
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1649977179
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1649977179
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1649977179
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_685
timestamp 1649977179
transform 1 0 64124 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_693
timestamp 1649977179
transform 1 0 64860 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_715
timestamp 1649977179
transform 1 0 66884 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1649977179
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1649977179
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1649977179
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1649977179
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1649977179
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1649977179
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1649977179
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1649977179
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1649977179
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_821
timestamp 1649977179
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1649977179
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1649977179
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_841
timestamp 1649977179
transform 1 0 78476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_853
timestamp 1649977179
transform 1 0 79580 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_865
timestamp 1649977179
transform 1 0 80684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_877
timestamp 1649977179
transform 1 0 81788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_889
timestamp 1649977179
transform 1 0 82892 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_895
timestamp 1649977179
transform 1 0 83444 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_897
timestamp 1649977179
transform 1 0 83628 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_909
timestamp 1649977179
transform 1 0 84732 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_921
timestamp 1649977179
transform 1 0 85836 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_933
timestamp 1649977179
transform 1 0 86940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_945
timestamp 1649977179
transform 1 0 88044 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_951
timestamp 1649977179
transform 1 0 88596 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_953
timestamp 1649977179
transform 1 0 88780 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_965
timestamp 1649977179
transform 1 0 89884 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_977
timestamp 1649977179
transform 1 0 90988 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_989
timestamp 1649977179
transform 1 0 92092 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1001
timestamp 1649977179
transform 1 0 93196 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1007
timestamp 1649977179
transform 1 0 93748 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1009
timestamp 1649977179
transform 1 0 93932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1021
timestamp 1649977179
transform 1 0 95036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1033
timestamp 1649977179
transform 1 0 96140 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1045
timestamp 1649977179
transform 1 0 97244 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1057
timestamp 1649977179
transform 1 0 98348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1063
timestamp 1649977179
transform 1 0 98900 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1065
timestamp 1649977179
transform 1 0 99084 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1077
timestamp 1649977179
transform 1 0 100188 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1089
timestamp 1649977179
transform 1 0 101292 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1101
timestamp 1649977179
transform 1 0 102396 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1113
timestamp 1649977179
transform 1 0 103500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1119
timestamp 1649977179
transform 1 0 104052 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1121
timestamp 1649977179
transform 1 0 104236 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1133
timestamp 1649977179
transform 1 0 105340 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1145
timestamp 1649977179
transform 1 0 106444 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1157
timestamp 1649977179
transform 1 0 107548 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1169
timestamp 1649977179
transform 1 0 108652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1175
timestamp 1649977179
transform 1 0 109204 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1177
timestamp 1649977179
transform 1 0 109388 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1189
timestamp 1649977179
transform 1 0 110492 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1201
timestamp 1649977179
transform 1 0 111596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1213
timestamp 1649977179
transform 1 0 112700 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1225
timestamp 1649977179
transform 1 0 113804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1231
timestamp 1649977179
transform 1 0 114356 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1233
timestamp 1649977179
transform 1 0 114540 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1245
timestamp 1649977179
transform 1 0 115644 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1257
timestamp 1649977179
transform 1 0 116748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1269
timestamp 1649977179
transform 1 0 117852 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_91
timestamp 1649977179
transform 1 0 9476 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_103
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_115
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_127
timestamp 1649977179
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1649977179
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_449
timestamp 1649977179
transform 1 0 42412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_460
timestamp 1649977179
transform 1 0 43424 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_472
timestamp 1649977179
transform 1 0 44528 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1649977179
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1649977179
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1649977179
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1649977179
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1649977179
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1649977179
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1649977179
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_725
timestamp 1649977179
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_737
timestamp 1649977179
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1649977179
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1649977179
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1649977179
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1649977179
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1649977179
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1649977179
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1649977179
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1649977179
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_813
timestamp 1649977179
transform 1 0 75900 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_825
timestamp 1649977179
transform 1 0 77004 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_837
timestamp 1649977179
transform 1 0 78108 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_849
timestamp 1649977179
transform 1 0 79212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_861
timestamp 1649977179
transform 1 0 80316 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_867
timestamp 1649977179
transform 1 0 80868 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_869
timestamp 1649977179
transform 1 0 81052 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_881
timestamp 1649977179
transform 1 0 82156 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_893
timestamp 1649977179
transform 1 0 83260 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_905
timestamp 1649977179
transform 1 0 84364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_917
timestamp 1649977179
transform 1 0 85468 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_923
timestamp 1649977179
transform 1 0 86020 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_925
timestamp 1649977179
transform 1 0 86204 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_937
timestamp 1649977179
transform 1 0 87308 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_949
timestamp 1649977179
transform 1 0 88412 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_961
timestamp 1649977179
transform 1 0 89516 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_973
timestamp 1649977179
transform 1 0 90620 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_979
timestamp 1649977179
transform 1 0 91172 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_981
timestamp 1649977179
transform 1 0 91356 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_993
timestamp 1649977179
transform 1 0 92460 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1005
timestamp 1649977179
transform 1 0 93564 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1017
timestamp 1649977179
transform 1 0 94668 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1029
timestamp 1649977179
transform 1 0 95772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1035
timestamp 1649977179
transform 1 0 96324 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1037
timestamp 1649977179
transform 1 0 96508 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1049
timestamp 1649977179
transform 1 0 97612 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1061
timestamp 1649977179
transform 1 0 98716 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1073
timestamp 1649977179
transform 1 0 99820 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1085
timestamp 1649977179
transform 1 0 100924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1091
timestamp 1649977179
transform 1 0 101476 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1093
timestamp 1649977179
transform 1 0 101660 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1105
timestamp 1649977179
transform 1 0 102764 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1117
timestamp 1649977179
transform 1 0 103868 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1129
timestamp 1649977179
transform 1 0 104972 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1141
timestamp 1649977179
transform 1 0 106076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1147
timestamp 1649977179
transform 1 0 106628 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1149
timestamp 1649977179
transform 1 0 106812 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1161
timestamp 1649977179
transform 1 0 107916 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1173
timestamp 1649977179
transform 1 0 109020 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1185
timestamp 1649977179
transform 1 0 110124 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1197
timestamp 1649977179
transform 1 0 111228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1203
timestamp 1649977179
transform 1 0 111780 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1205
timestamp 1649977179
transform 1 0 111964 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1217
timestamp 1649977179
transform 1 0 113068 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1229
timestamp 1649977179
transform 1 0 114172 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1241
timestamp 1649977179
transform 1 0 115276 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1253
timestamp 1649977179
transform 1 0 116380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1259
timestamp 1649977179
transform 1 0 116932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1261
timestamp 1649977179
transform 1 0 117116 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1269
timestamp 1649977179
transform 1 0 117852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1273
timestamp 1649977179
transform 1 0 118220 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_6
timestamp 1649977179
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_18
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_30
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_42
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_408
timestamp 1649977179
transform 1 0 38640 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_419
timestamp 1649977179
transform 1 0 39652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1649977179
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1649977179
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1649977179
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1649977179
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1649977179
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1649977179
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1649977179
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1649977179
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1649977179
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1649977179
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_729
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_741
timestamp 1649977179
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_753
timestamp 1649977179
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_765
timestamp 1649977179
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1649977179
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1649977179
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1649977179
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1649977179
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_809
timestamp 1649977179
transform 1 0 75532 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_821
timestamp 1649977179
transform 1 0 76636 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_827
timestamp 1649977179
transform 1 0 77188 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_839
timestamp 1649977179
transform 1 0 78292 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_841
timestamp 1649977179
transform 1 0 78476 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_853
timestamp 1649977179
transform 1 0 79580 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_865
timestamp 1649977179
transform 1 0 80684 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_877
timestamp 1649977179
transform 1 0 81788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_889
timestamp 1649977179
transform 1 0 82892 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_895
timestamp 1649977179
transform 1 0 83444 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_897
timestamp 1649977179
transform 1 0 83628 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_909
timestamp 1649977179
transform 1 0 84732 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_921
timestamp 1649977179
transform 1 0 85836 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_933
timestamp 1649977179
transform 1 0 86940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_945
timestamp 1649977179
transform 1 0 88044 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_951
timestamp 1649977179
transform 1 0 88596 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_953
timestamp 1649977179
transform 1 0 88780 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_965
timestamp 1649977179
transform 1 0 89884 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_977
timestamp 1649977179
transform 1 0 90988 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_989
timestamp 1649977179
transform 1 0 92092 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1001
timestamp 1649977179
transform 1 0 93196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1007
timestamp 1649977179
transform 1 0 93748 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1009
timestamp 1649977179
transform 1 0 93932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1021
timestamp 1649977179
transform 1 0 95036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1033
timestamp 1649977179
transform 1 0 96140 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1045
timestamp 1649977179
transform 1 0 97244 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1057
timestamp 1649977179
transform 1 0 98348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1063
timestamp 1649977179
transform 1 0 98900 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1065
timestamp 1649977179
transform 1 0 99084 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1077
timestamp 1649977179
transform 1 0 100188 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1089
timestamp 1649977179
transform 1 0 101292 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1101
timestamp 1649977179
transform 1 0 102396 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1113
timestamp 1649977179
transform 1 0 103500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1119
timestamp 1649977179
transform 1 0 104052 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1121
timestamp 1649977179
transform 1 0 104236 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1133
timestamp 1649977179
transform 1 0 105340 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1145
timestamp 1649977179
transform 1 0 106444 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1157
timestamp 1649977179
transform 1 0 107548 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1169
timestamp 1649977179
transform 1 0 108652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1175
timestamp 1649977179
transform 1 0 109204 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1177
timestamp 1649977179
transform 1 0 109388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1189
timestamp 1649977179
transform 1 0 110492 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1201
timestamp 1649977179
transform 1 0 111596 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1213
timestamp 1649977179
transform 1 0 112700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1225
timestamp 1649977179
transform 1 0 113804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1231
timestamp 1649977179
transform 1 0 114356 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1233
timestamp 1649977179
transform 1 0 114540 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1245
timestamp 1649977179
transform 1 0 115644 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1257
timestamp 1649977179
transform 1 0 116748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1273
timestamp 1649977179
transform 1 0 118220 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1649977179
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_237
timestamp 1649977179
transform 1 0 22908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1649977179
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_325
timestamp 1649977179
transform 1 0 31004 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_336
timestamp 1649977179
transform 1 0 32016 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_348
timestamp 1649977179
transform 1 0 33120 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1649977179
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1649977179
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1649977179
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1649977179
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1649977179
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1649977179
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1649977179
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1649977179
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1649977179
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_713
timestamp 1649977179
transform 1 0 66700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_722
timestamp 1649977179
transform 1 0 67528 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_726
timestamp 1649977179
transform 1 0 67896 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_732
timestamp 1649977179
transform 1 0 68448 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_744
timestamp 1649977179
transform 1 0 69552 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_757
timestamp 1649977179
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_769
timestamp 1649977179
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_781
timestamp 1649977179
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_793
timestamp 1649977179
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 1649977179
transform 1 0 75164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 1649977179
transform 1 0 75716 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_813
timestamp 1649977179
transform 1 0 75900 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_825
timestamp 1649977179
transform 1 0 77004 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_837
timestamp 1649977179
transform 1 0 78108 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_849
timestamp 1649977179
transform 1 0 79212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_861
timestamp 1649977179
transform 1 0 80316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_867
timestamp 1649977179
transform 1 0 80868 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_869
timestamp 1649977179
transform 1 0 81052 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_881
timestamp 1649977179
transform 1 0 82156 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_893
timestamp 1649977179
transform 1 0 83260 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_905
timestamp 1649977179
transform 1 0 84364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_917
timestamp 1649977179
transform 1 0 85468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_923
timestamp 1649977179
transform 1 0 86020 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_925
timestamp 1649977179
transform 1 0 86204 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_937
timestamp 1649977179
transform 1 0 87308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_949
timestamp 1649977179
transform 1 0 88412 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_961
timestamp 1649977179
transform 1 0 89516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_973
timestamp 1649977179
transform 1 0 90620 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_979
timestamp 1649977179
transform 1 0 91172 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_981
timestamp 1649977179
transform 1 0 91356 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_993
timestamp 1649977179
transform 1 0 92460 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1005
timestamp 1649977179
transform 1 0 93564 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1017
timestamp 1649977179
transform 1 0 94668 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1029
timestamp 1649977179
transform 1 0 95772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1035
timestamp 1649977179
transform 1 0 96324 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1037
timestamp 1649977179
transform 1 0 96508 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1049
timestamp 1649977179
transform 1 0 97612 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1061
timestamp 1649977179
transform 1 0 98716 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1073
timestamp 1649977179
transform 1 0 99820 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1085
timestamp 1649977179
transform 1 0 100924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1091
timestamp 1649977179
transform 1 0 101476 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1093
timestamp 1649977179
transform 1 0 101660 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1105
timestamp 1649977179
transform 1 0 102764 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1117
timestamp 1649977179
transform 1 0 103868 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1129
timestamp 1649977179
transform 1 0 104972 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1141
timestamp 1649977179
transform 1 0 106076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1147
timestamp 1649977179
transform 1 0 106628 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1149
timestamp 1649977179
transform 1 0 106812 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1161
timestamp 1649977179
transform 1 0 107916 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1173
timestamp 1649977179
transform 1 0 109020 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1185
timestamp 1649977179
transform 1 0 110124 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1197
timestamp 1649977179
transform 1 0 111228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1203
timestamp 1649977179
transform 1 0 111780 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1205
timestamp 1649977179
transform 1 0 111964 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1217
timestamp 1649977179
transform 1 0 113068 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1229
timestamp 1649977179
transform 1 0 114172 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1241
timestamp 1649977179
transform 1 0 115276 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1253
timestamp 1649977179
transform 1 0 116380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1259
timestamp 1649977179
transform 1 0 116932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1261
timestamp 1649977179
transform 1 0 117116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1273
timestamp 1649977179
transform 1 0 118220 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_6
timestamp 1649977179
transform 1 0 1656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_18
timestamp 1649977179
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_30
timestamp 1649977179
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_42
timestamp 1649977179
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_340
timestamp 1649977179
transform 1 0 32384 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_352
timestamp 1649977179
transform 1 0 33488 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_364
timestamp 1649977179
transform 1 0 34592 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_376
timestamp 1649977179
transform 1 0 35696 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1649977179
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1649977179
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1649977179
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1649977179
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1649977179
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1649977179
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_697
timestamp 1649977179
transform 1 0 65228 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_705
timestamp 1649977179
transform 1 0 65964 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_724
timestamp 1649977179
transform 1 0 67712 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_736
timestamp 1649977179
transform 1 0 68816 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_742
timestamp 1649977179
transform 1 0 69368 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_749
timestamp 1649977179
transform 1 0 70012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_761
timestamp 1649977179
transform 1 0 71116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_773
timestamp 1649977179
transform 1 0 72220 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_781
timestamp 1649977179
transform 1 0 72956 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1649977179
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_797
timestamp 1649977179
transform 1 0 74428 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_809
timestamp 1649977179
transform 1 0 75532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_813
timestamp 1649977179
transform 1 0 75900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_816
timestamp 1649977179
transform 1 0 76176 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_827
timestamp 1649977179
transform 1 0 77188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_839
timestamp 1649977179
transform 1 0 78292 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_841
timestamp 1649977179
transform 1 0 78476 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_853
timestamp 1649977179
transform 1 0 79580 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_865
timestamp 1649977179
transform 1 0 80684 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_877
timestamp 1649977179
transform 1 0 81788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_889
timestamp 1649977179
transform 1 0 82892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_895
timestamp 1649977179
transform 1 0 83444 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_897
timestamp 1649977179
transform 1 0 83628 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_909
timestamp 1649977179
transform 1 0 84732 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_921
timestamp 1649977179
transform 1 0 85836 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_933
timestamp 1649977179
transform 1 0 86940 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_945
timestamp 1649977179
transform 1 0 88044 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_951
timestamp 1649977179
transform 1 0 88596 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_953
timestamp 1649977179
transform 1 0 88780 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_965
timestamp 1649977179
transform 1 0 89884 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_977
timestamp 1649977179
transform 1 0 90988 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_989
timestamp 1649977179
transform 1 0 92092 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1001
timestamp 1649977179
transform 1 0 93196 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1007
timestamp 1649977179
transform 1 0 93748 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1009
timestamp 1649977179
transform 1 0 93932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1021
timestamp 1649977179
transform 1 0 95036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1033
timestamp 1649977179
transform 1 0 96140 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1045
timestamp 1649977179
transform 1 0 97244 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1057
timestamp 1649977179
transform 1 0 98348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1063
timestamp 1649977179
transform 1 0 98900 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1065
timestamp 1649977179
transform 1 0 99084 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1077
timestamp 1649977179
transform 1 0 100188 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1089
timestamp 1649977179
transform 1 0 101292 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1101
timestamp 1649977179
transform 1 0 102396 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1113
timestamp 1649977179
transform 1 0 103500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1119
timestamp 1649977179
transform 1 0 104052 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1121
timestamp 1649977179
transform 1 0 104236 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1133
timestamp 1649977179
transform 1 0 105340 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1145
timestamp 1649977179
transform 1 0 106444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1157
timestamp 1649977179
transform 1 0 107548 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1161
timestamp 1649977179
transform 1 0 107916 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1165
timestamp 1649977179
transform 1 0 108284 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1173
timestamp 1649977179
transform 1 0 109020 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1177
timestamp 1649977179
transform 1 0 109388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1189
timestamp 1649977179
transform 1 0 110492 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1201
timestamp 1649977179
transform 1 0 111596 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1213
timestamp 1649977179
transform 1 0 112700 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1225
timestamp 1649977179
transform 1 0 113804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1231
timestamp 1649977179
transform 1 0 114356 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1233
timestamp 1649977179
transform 1 0 114540 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1245
timestamp 1649977179
transform 1 0 115644 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1257
timestamp 1649977179
transform 1 0 116748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1269
timestamp 1649977179
transform 1 0 117852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1649977179
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1649977179
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1649977179
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1649977179
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1649977179
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1649977179
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1649977179
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1649977179
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1649977179
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1649977179
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_713
timestamp 1649977179
transform 1 0 66700 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_721
timestamp 1649977179
transform 1 0 67436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_743
timestamp 1649977179
transform 1 0 69460 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_752
timestamp 1649977179
transform 1 0 70288 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_757
timestamp 1649977179
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_769
timestamp 1649977179
transform 1 0 71852 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_781
timestamp 1649977179
transform 1 0 72956 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_793
timestamp 1649977179
transform 1 0 74060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 1649977179
transform 1 0 75164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 1649977179
transform 1 0 75716 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_813
timestamp 1649977179
transform 1 0 75900 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_825
timestamp 1649977179
transform 1 0 77004 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_837
timestamp 1649977179
transform 1 0 78108 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_849
timestamp 1649977179
transform 1 0 79212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_861
timestamp 1649977179
transform 1 0 80316 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_867
timestamp 1649977179
transform 1 0 80868 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_869
timestamp 1649977179
transform 1 0 81052 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_881
timestamp 1649977179
transform 1 0 82156 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_893
timestamp 1649977179
transform 1 0 83260 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_905
timestamp 1649977179
transform 1 0 84364 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_917
timestamp 1649977179
transform 1 0 85468 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_923
timestamp 1649977179
transform 1 0 86020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_925
timestamp 1649977179
transform 1 0 86204 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_932
timestamp 1649977179
transform 1 0 86848 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_944
timestamp 1649977179
transform 1 0 87952 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_956
timestamp 1649977179
transform 1 0 89056 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_968
timestamp 1649977179
transform 1 0 90160 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_981
timestamp 1649977179
transform 1 0 91356 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_993
timestamp 1649977179
transform 1 0 92460 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1005
timestamp 1649977179
transform 1 0 93564 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1017
timestamp 1649977179
transform 1 0 94668 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1029
timestamp 1649977179
transform 1 0 95772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1035
timestamp 1649977179
transform 1 0 96324 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1037
timestamp 1649977179
transform 1 0 96508 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1049
timestamp 1649977179
transform 1 0 97612 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1061
timestamp 1649977179
transform 1 0 98716 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1073
timestamp 1649977179
transform 1 0 99820 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1085
timestamp 1649977179
transform 1 0 100924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1091
timestamp 1649977179
transform 1 0 101476 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1093
timestamp 1649977179
transform 1 0 101660 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1105
timestamp 1649977179
transform 1 0 102764 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1117
timestamp 1649977179
transform 1 0 103868 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1129
timestamp 1649977179
transform 1 0 104972 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1141
timestamp 1649977179
transform 1 0 106076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1147
timestamp 1649977179
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1149
timestamp 1649977179
transform 1 0 106812 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1161
timestamp 1649977179
transform 1 0 107916 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1173
timestamp 1649977179
transform 1 0 109020 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1185
timestamp 1649977179
transform 1 0 110124 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1197
timestamp 1649977179
transform 1 0 111228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1203
timestamp 1649977179
transform 1 0 111780 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1205
timestamp 1649977179
transform 1 0 111964 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1217
timestamp 1649977179
transform 1 0 113068 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1229
timestamp 1649977179
transform 1 0 114172 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1241
timestamp 1649977179
transform 1 0 115276 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1253
timestamp 1649977179
transform 1 0 116380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1259
timestamp 1649977179
transform 1 0 116932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1261
timestamp 1649977179
transform 1 0 117116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1269
timestamp 1649977179
transform 1 0 117852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1273
timestamp 1649977179
transform 1 0 118220 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1649977179
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1649977179
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1649977179
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1649977179
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1649977179
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1649977179
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1649977179
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_697
timestamp 1649977179
transform 1 0 65228 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_704
timestamp 1649977179
transform 1 0 65872 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_724
timestamp 1649977179
transform 1 0 67712 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1649977179
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_753
timestamp 1649977179
transform 1 0 70380 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_763
timestamp 1649977179
transform 1 0 71300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_775
timestamp 1649977179
transform 1 0 72404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 1649977179
transform 1 0 73140 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_785
timestamp 1649977179
transform 1 0 73324 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_797
timestamp 1649977179
transform 1 0 74428 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_809
timestamp 1649977179
transform 1 0 75532 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_821
timestamp 1649977179
transform 1 0 76636 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_833
timestamp 1649977179
transform 1 0 77740 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_839
timestamp 1649977179
transform 1 0 78292 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_841
timestamp 1649977179
transform 1 0 78476 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_853
timestamp 1649977179
transform 1 0 79580 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_865
timestamp 1649977179
transform 1 0 80684 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_877
timestamp 1649977179
transform 1 0 81788 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_889
timestamp 1649977179
transform 1 0 82892 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_895
timestamp 1649977179
transform 1 0 83444 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_897
timestamp 1649977179
transform 1 0 83628 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_909
timestamp 1649977179
transform 1 0 84732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_919
timestamp 1649977179
transform 1 0 85652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_930
timestamp 1649977179
transform 1 0 86664 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_942
timestamp 1649977179
transform 1 0 87768 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_950
timestamp 1649977179
transform 1 0 88504 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_953
timestamp 1649977179
transform 1 0 88780 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_965
timestamp 1649977179
transform 1 0 89884 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_977
timestamp 1649977179
transform 1 0 90988 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_989
timestamp 1649977179
transform 1 0 92092 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1001
timestamp 1649977179
transform 1 0 93196 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1007
timestamp 1649977179
transform 1 0 93748 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1009
timestamp 1649977179
transform 1 0 93932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1021
timestamp 1649977179
transform 1 0 95036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1033
timestamp 1649977179
transform 1 0 96140 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1045
timestamp 1649977179
transform 1 0 97244 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1057
timestamp 1649977179
transform 1 0 98348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1063
timestamp 1649977179
transform 1 0 98900 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1065
timestamp 1649977179
transform 1 0 99084 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1077
timestamp 1649977179
transform 1 0 100188 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1089
timestamp 1649977179
transform 1 0 101292 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1101
timestamp 1649977179
transform 1 0 102396 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1113
timestamp 1649977179
transform 1 0 103500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1119
timestamp 1649977179
transform 1 0 104052 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1121
timestamp 1649977179
transform 1 0 104236 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1133
timestamp 1649977179
transform 1 0 105340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1145
timestamp 1649977179
transform 1 0 106444 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1151
timestamp 1649977179
transform 1 0 106996 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1156
timestamp 1649977179
transform 1 0 107456 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1168
timestamp 1649977179
transform 1 0 108560 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1177
timestamp 1649977179
transform 1 0 109388 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1189
timestamp 1649977179
transform 1 0 110492 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1201
timestamp 1649977179
transform 1 0 111596 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1213
timestamp 1649977179
transform 1 0 112700 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1225
timestamp 1649977179
transform 1 0 113804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1231
timestamp 1649977179
transform 1 0 114356 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1233
timestamp 1649977179
transform 1 0 114540 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1245
timestamp 1649977179
transform 1 0 115644 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1257
timestamp 1649977179
transform 1 0 116748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_1273
timestamp 1649977179
transform 1 0 118220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_6
timestamp 1649977179
transform 1 0 1656 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_543
timestamp 1649977179
transform 1 0 51060 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_555
timestamp 1649977179
transform 1 0 52164 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_567
timestamp 1649977179
transform 1 0 53268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_579
timestamp 1649977179
transform 1 0 54372 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_593
timestamp 1649977179
transform 1 0 55660 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_605
timestamp 1649977179
transform 1 0 56764 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_617
timestamp 1649977179
transform 1 0 57868 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_629
timestamp 1649977179
transform 1 0 58972 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_641
timestamp 1649977179
transform 1 0 60076 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1649977179
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1649977179
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1649977179
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_681
timestamp 1649977179
transform 1 0 63756 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_689
timestamp 1649977179
transform 1 0 64492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_696
timestamp 1649977179
transform 1 0 65136 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_701
timestamp 1649977179
transform 1 0 65596 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_710
timestamp 1649977179
transform 1 0 66424 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_730
timestamp 1649977179
transform 1 0 68264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_750
timestamp 1649977179
transform 1 0 70104 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_761
timestamp 1649977179
transform 1 0 71116 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_768
timestamp 1649977179
transform 1 0 71760 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_780
timestamp 1649977179
transform 1 0 72864 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_792
timestamp 1649977179
transform 1 0 73968 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_804
timestamp 1649977179
transform 1 0 75072 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_813
timestamp 1649977179
transform 1 0 75900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_825
timestamp 1649977179
transform 1 0 77004 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_837
timestamp 1649977179
transform 1 0 78108 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_849
timestamp 1649977179
transform 1 0 79212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_861
timestamp 1649977179
transform 1 0 80316 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_867
timestamp 1649977179
transform 1 0 80868 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_869
timestamp 1649977179
transform 1 0 81052 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_881
timestamp 1649977179
transform 1 0 82156 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_893
timestamp 1649977179
transform 1 0 83260 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_905
timestamp 1649977179
transform 1 0 84364 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_917
timestamp 1649977179
transform 1 0 85468 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_923
timestamp 1649977179
transform 1 0 86020 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_925
timestamp 1649977179
transform 1 0 86204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_937
timestamp 1649977179
transform 1 0 87308 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_949
timestamp 1649977179
transform 1 0 88412 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_961
timestamp 1649977179
transform 1 0 89516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_973
timestamp 1649977179
transform 1 0 90620 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_979
timestamp 1649977179
transform 1 0 91172 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_981
timestamp 1649977179
transform 1 0 91356 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_993
timestamp 1649977179
transform 1 0 92460 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1005
timestamp 1649977179
transform 1 0 93564 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1017
timestamp 1649977179
transform 1 0 94668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1029
timestamp 1649977179
transform 1 0 95772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1035
timestamp 1649977179
transform 1 0 96324 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1037
timestamp 1649977179
transform 1 0 96508 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1049
timestamp 1649977179
transform 1 0 97612 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1061
timestamp 1649977179
transform 1 0 98716 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1073
timestamp 1649977179
transform 1 0 99820 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1085
timestamp 1649977179
transform 1 0 100924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1091
timestamp 1649977179
transform 1 0 101476 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1093
timestamp 1649977179
transform 1 0 101660 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1105
timestamp 1649977179
transform 1 0 102764 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1117
timestamp 1649977179
transform 1 0 103868 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1129
timestamp 1649977179
transform 1 0 104972 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1141
timestamp 1649977179
transform 1 0 106076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1147
timestamp 1649977179
transform 1 0 106628 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1149
timestamp 1649977179
transform 1 0 106812 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1161
timestamp 1649977179
transform 1 0 107916 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1173
timestamp 1649977179
transform 1 0 109020 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1185
timestamp 1649977179
transform 1 0 110124 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1197
timestamp 1649977179
transform 1 0 111228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1203
timestamp 1649977179
transform 1 0 111780 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1205
timestamp 1649977179
transform 1 0 111964 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1217
timestamp 1649977179
transform 1 0 113068 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1229
timestamp 1649977179
transform 1 0 114172 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1241
timestamp 1649977179
transform 1 0 115276 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1253
timestamp 1649977179
transform 1 0 116380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1259
timestamp 1649977179
transform 1 0 116932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_1261
timestamp 1649977179
transform 1 0 117116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_1273
timestamp 1649977179
transform 1 0 118220 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_78
timestamp 1649977179
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_90
timestamp 1649977179
transform 1 0 9384 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_525
timestamp 1649977179
transform 1 0 49404 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_532
timestamp 1649977179
transform 1 0 50048 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_542
timestamp 1649977179
transform 1 0 50968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_554
timestamp 1649977179
transform 1 0 52072 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_569
timestamp 1649977179
transform 1 0 53452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_577
timestamp 1649977179
transform 1 0 54188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_591
timestamp 1649977179
transform 1 0 55476 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_601
timestamp 1649977179
transform 1 0 56396 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_613
timestamp 1649977179
transform 1 0 57500 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1649977179
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1649977179
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1649977179
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1649977179
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1649977179
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_673
timestamp 1649977179
transform 1 0 63020 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_681
timestamp 1649977179
transform 1 0 63756 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_689
timestamp 1649977179
transform 1 0 64492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_699
timestamp 1649977179
transform 1 0 65412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_709
timestamp 1649977179
transform 1 0 66332 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_713
timestamp 1649977179
transform 1 0 66700 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_724
timestamp 1649977179
transform 1 0 67712 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1649977179
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_733
timestamp 1649977179
transform 1 0 68540 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_744
timestamp 1649977179
transform 1 0 69552 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_753
timestamp 1649977179
transform 1 0 70380 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_760
timestamp 1649977179
transform 1 0 71024 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_772
timestamp 1649977179
transform 1 0 72128 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_785
timestamp 1649977179
transform 1 0 73324 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_797
timestamp 1649977179
transform 1 0 74428 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_809
timestamp 1649977179
transform 1 0 75532 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_821
timestamp 1649977179
transform 1 0 76636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_833
timestamp 1649977179
transform 1 0 77740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_839
timestamp 1649977179
transform 1 0 78292 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_841
timestamp 1649977179
transform 1 0 78476 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_853
timestamp 1649977179
transform 1 0 79580 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_865
timestamp 1649977179
transform 1 0 80684 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_877
timestamp 1649977179
transform 1 0 81788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_889
timestamp 1649977179
transform 1 0 82892 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_895
timestamp 1649977179
transform 1 0 83444 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_897
timestamp 1649977179
transform 1 0 83628 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_909
timestamp 1649977179
transform 1 0 84732 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_921
timestamp 1649977179
transform 1 0 85836 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_933
timestamp 1649977179
transform 1 0 86940 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_945
timestamp 1649977179
transform 1 0 88044 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_951
timestamp 1649977179
transform 1 0 88596 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_953
timestamp 1649977179
transform 1 0 88780 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_965
timestamp 1649977179
transform 1 0 89884 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_977
timestamp 1649977179
transform 1 0 90988 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_989
timestamp 1649977179
transform 1 0 92092 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1001
timestamp 1649977179
transform 1 0 93196 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1007
timestamp 1649977179
transform 1 0 93748 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1009
timestamp 1649977179
transform 1 0 93932 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1021
timestamp 1649977179
transform 1 0 95036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1033
timestamp 1649977179
transform 1 0 96140 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1045
timestamp 1649977179
transform 1 0 97244 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1057
timestamp 1649977179
transform 1 0 98348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1063
timestamp 1649977179
transform 1 0 98900 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1065
timestamp 1649977179
transform 1 0 99084 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1077
timestamp 1649977179
transform 1 0 100188 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1089
timestamp 1649977179
transform 1 0 101292 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1101
timestamp 1649977179
transform 1 0 102396 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1113
timestamp 1649977179
transform 1 0 103500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1119
timestamp 1649977179
transform 1 0 104052 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1121
timestamp 1649977179
transform 1 0 104236 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1133
timestamp 1649977179
transform 1 0 105340 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1145
timestamp 1649977179
transform 1 0 106444 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1157
timestamp 1649977179
transform 1 0 107548 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1169
timestamp 1649977179
transform 1 0 108652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1175
timestamp 1649977179
transform 1 0 109204 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1177
timestamp 1649977179
transform 1 0 109388 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1189
timestamp 1649977179
transform 1 0 110492 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1201
timestamp 1649977179
transform 1 0 111596 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1213
timestamp 1649977179
transform 1 0 112700 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1225
timestamp 1649977179
transform 1 0 113804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1231
timestamp 1649977179
transform 1 0 114356 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1233
timestamp 1649977179
transform 1 0 114540 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1245
timestamp 1649977179
transform 1 0 115644 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1257
timestamp 1649977179
transform 1 0 116748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_1269
timestamp 1649977179
transform 1 0 117852 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_6
timestamp 1649977179
transform 1 0 1656 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1649977179
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_317
timestamp 1649977179
transform 1 0 30268 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_324
timestamp 1649977179
transform 1 0 30912 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_336
timestamp 1649977179
transform 1 0 32016 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_348
timestamp 1649977179
transform 1 0 33120 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1649977179
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1649977179
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1649977179
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1649977179
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1649977179
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1649977179
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1649977179
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_681
timestamp 1649977179
transform 1 0 63756 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_689
timestamp 1649977179
transform 1 0 64492 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_694
timestamp 1649977179
transform 1 0 64952 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_710
timestamp 1649977179
transform 1 0 66424 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_714
timestamp 1649977179
transform 1 0 66792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_723
timestamp 1649977179
transform 1 0 67620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_734
timestamp 1649977179
transform 1 0 68632 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_738
timestamp 1649977179
transform 1 0 69000 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_745
timestamp 1649977179
transform 1 0 69644 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_753
timestamp 1649977179
transform 1 0 70380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_766
timestamp 1649977179
transform 1 0 71576 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_770
timestamp 1649977179
transform 1 0 71944 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_782
timestamp 1649977179
transform 1 0 73048 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_794
timestamp 1649977179
transform 1 0 74152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_806
timestamp 1649977179
transform 1 0 75256 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_813
timestamp 1649977179
transform 1 0 75900 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_825
timestamp 1649977179
transform 1 0 77004 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_837
timestamp 1649977179
transform 1 0 78108 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_849
timestamp 1649977179
transform 1 0 79212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_861
timestamp 1649977179
transform 1 0 80316 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_867
timestamp 1649977179
transform 1 0 80868 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_869
timestamp 1649977179
transform 1 0 81052 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_881
timestamp 1649977179
transform 1 0 82156 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_893
timestamp 1649977179
transform 1 0 83260 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_905
timestamp 1649977179
transform 1 0 84364 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_917
timestamp 1649977179
transform 1 0 85468 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_923
timestamp 1649977179
transform 1 0 86020 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_925
timestamp 1649977179
transform 1 0 86204 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_937
timestamp 1649977179
transform 1 0 87308 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_949
timestamp 1649977179
transform 1 0 88412 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_961
timestamp 1649977179
transform 1 0 89516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_973
timestamp 1649977179
transform 1 0 90620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_979
timestamp 1649977179
transform 1 0 91172 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_981
timestamp 1649977179
transform 1 0 91356 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_993
timestamp 1649977179
transform 1 0 92460 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1005
timestamp 1649977179
transform 1 0 93564 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1017
timestamp 1649977179
transform 1 0 94668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1029
timestamp 1649977179
transform 1 0 95772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1035
timestamp 1649977179
transform 1 0 96324 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1037
timestamp 1649977179
transform 1 0 96508 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1049
timestamp 1649977179
transform 1 0 97612 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1061
timestamp 1649977179
transform 1 0 98716 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1073
timestamp 1649977179
transform 1 0 99820 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1085
timestamp 1649977179
transform 1 0 100924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1091
timestamp 1649977179
transform 1 0 101476 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1093
timestamp 1649977179
transform 1 0 101660 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1105
timestamp 1649977179
transform 1 0 102764 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1117
timestamp 1649977179
transform 1 0 103868 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1129
timestamp 1649977179
transform 1 0 104972 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1141
timestamp 1649977179
transform 1 0 106076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1147
timestamp 1649977179
transform 1 0 106628 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1149
timestamp 1649977179
transform 1 0 106812 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1161
timestamp 1649977179
transform 1 0 107916 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1173
timestamp 1649977179
transform 1 0 109020 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1185
timestamp 1649977179
transform 1 0 110124 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1197
timestamp 1649977179
transform 1 0 111228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1203
timestamp 1649977179
transform 1 0 111780 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1205
timestamp 1649977179
transform 1 0 111964 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1217
timestamp 1649977179
transform 1 0 113068 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1229
timestamp 1649977179
transform 1 0 114172 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1241
timestamp 1649977179
transform 1 0 115276 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1253
timestamp 1649977179
transform 1 0 116380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1259
timestamp 1649977179
transform 1 0 116932 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1261
timestamp 1649977179
transform 1 0 117116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_1273
timestamp 1649977179
transform 1 0 118220 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1649977179
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1649977179
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1649977179
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1649977179
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1649977179
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1649977179
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1649977179
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1649977179
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_709
timestamp 1649977179
transform 1 0 66332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_713
timestamp 1649977179
transform 1 0 66700 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_717
timestamp 1649977179
transform 1 0 67068 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_725
timestamp 1649977179
transform 1 0 67804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_734
timestamp 1649977179
transform 1 0 68632 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_740
timestamp 1649977179
transform 1 0 69184 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_745
timestamp 1649977179
transform 1 0 69644 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_757
timestamp 1649977179
transform 1 0 70748 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_769
timestamp 1649977179
transform 1 0 71852 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_781
timestamp 1649977179
transform 1 0 72956 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_785
timestamp 1649977179
transform 1 0 73324 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_797
timestamp 1649977179
transform 1 0 74428 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_809
timestamp 1649977179
transform 1 0 75532 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_821
timestamp 1649977179
transform 1 0 76636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_833
timestamp 1649977179
transform 1 0 77740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_839
timestamp 1649977179
transform 1 0 78292 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_841
timestamp 1649977179
transform 1 0 78476 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_853
timestamp 1649977179
transform 1 0 79580 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_865
timestamp 1649977179
transform 1 0 80684 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_877
timestamp 1649977179
transform 1 0 81788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_889
timestamp 1649977179
transform 1 0 82892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_895
timestamp 1649977179
transform 1 0 83444 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_897
timestamp 1649977179
transform 1 0 83628 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_909
timestamp 1649977179
transform 1 0 84732 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_921
timestamp 1649977179
transform 1 0 85836 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_933
timestamp 1649977179
transform 1 0 86940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_945
timestamp 1649977179
transform 1 0 88044 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_951
timestamp 1649977179
transform 1 0 88596 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_953
timestamp 1649977179
transform 1 0 88780 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_965
timestamp 1649977179
transform 1 0 89884 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_977
timestamp 1649977179
transform 1 0 90988 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_989
timestamp 1649977179
transform 1 0 92092 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1001
timestamp 1649977179
transform 1 0 93196 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1007
timestamp 1649977179
transform 1 0 93748 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1009
timestamp 1649977179
transform 1 0 93932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1021
timestamp 1649977179
transform 1 0 95036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1033
timestamp 1649977179
transform 1 0 96140 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1045
timestamp 1649977179
transform 1 0 97244 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1057
timestamp 1649977179
transform 1 0 98348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1063
timestamp 1649977179
transform 1 0 98900 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1065
timestamp 1649977179
transform 1 0 99084 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1077
timestamp 1649977179
transform 1 0 100188 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1089
timestamp 1649977179
transform 1 0 101292 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1101
timestamp 1649977179
transform 1 0 102396 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1113
timestamp 1649977179
transform 1 0 103500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1119
timestamp 1649977179
transform 1 0 104052 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1121
timestamp 1649977179
transform 1 0 104236 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1133
timestamp 1649977179
transform 1 0 105340 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1145
timestamp 1649977179
transform 1 0 106444 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1157
timestamp 1649977179
transform 1 0 107548 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1169
timestamp 1649977179
transform 1 0 108652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1175
timestamp 1649977179
transform 1 0 109204 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1177
timestamp 1649977179
transform 1 0 109388 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1189
timestamp 1649977179
transform 1 0 110492 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1201
timestamp 1649977179
transform 1 0 111596 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1213
timestamp 1649977179
transform 1 0 112700 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1225
timestamp 1649977179
transform 1 0 113804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1231
timestamp 1649977179
transform 1 0 114356 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1233
timestamp 1649977179
transform 1 0 114540 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1245
timestamp 1649977179
transform 1 0 115644 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1257
timestamp 1649977179
transform 1 0 116748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1269
timestamp 1649977179
transform 1 0 117852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_1273
timestamp 1649977179
transform 1 0 118220 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_6
timestamp 1649977179
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1649977179
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1649977179
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1649977179
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1649977179
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1649977179
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1649977179
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1649977179
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1649977179
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1649977179
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1649977179
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1649977179
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_713
timestamp 1649977179
transform 1 0 66700 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_719
timestamp 1649977179
transform 1 0 67252 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_731
timestamp 1649977179
transform 1 0 68356 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_743
timestamp 1649977179
transform 1 0 69460 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 1649977179
transform 1 0 70564 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_757
timestamp 1649977179
transform 1 0 70748 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_767
timestamp 1649977179
transform 1 0 71668 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_779
timestamp 1649977179
transform 1 0 72772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_791
timestamp 1649977179
transform 1 0 73876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_803
timestamp 1649977179
transform 1 0 74980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 1649977179
transform 1 0 75716 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_813
timestamp 1649977179
transform 1 0 75900 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_825
timestamp 1649977179
transform 1 0 77004 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_837
timestamp 1649977179
transform 1 0 78108 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_849
timestamp 1649977179
transform 1 0 79212 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_861
timestamp 1649977179
transform 1 0 80316 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_867
timestamp 1649977179
transform 1 0 80868 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_869
timestamp 1649977179
transform 1 0 81052 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_879
timestamp 1649977179
transform 1 0 81972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_890
timestamp 1649977179
transform 1 0 82984 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_894
timestamp 1649977179
transform 1 0 83352 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_906
timestamp 1649977179
transform 1 0 84456 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_918
timestamp 1649977179
transform 1 0 85560 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_925
timestamp 1649977179
transform 1 0 86204 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_937
timestamp 1649977179
transform 1 0 87308 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_949
timestamp 1649977179
transform 1 0 88412 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_961
timestamp 1649977179
transform 1 0 89516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_973
timestamp 1649977179
transform 1 0 90620 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_979
timestamp 1649977179
transform 1 0 91172 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_981
timestamp 1649977179
transform 1 0 91356 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_993
timestamp 1649977179
transform 1 0 92460 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1005
timestamp 1649977179
transform 1 0 93564 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1017
timestamp 1649977179
transform 1 0 94668 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1029
timestamp 1649977179
transform 1 0 95772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1035
timestamp 1649977179
transform 1 0 96324 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1037
timestamp 1649977179
transform 1 0 96508 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1049
timestamp 1649977179
transform 1 0 97612 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1061
timestamp 1649977179
transform 1 0 98716 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1073
timestamp 1649977179
transform 1 0 99820 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1085
timestamp 1649977179
transform 1 0 100924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1091
timestamp 1649977179
transform 1 0 101476 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1093
timestamp 1649977179
transform 1 0 101660 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1105
timestamp 1649977179
transform 1 0 102764 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1117
timestamp 1649977179
transform 1 0 103868 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1129
timestamp 1649977179
transform 1 0 104972 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1141
timestamp 1649977179
transform 1 0 106076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1147
timestamp 1649977179
transform 1 0 106628 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1149
timestamp 1649977179
transform 1 0 106812 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1161
timestamp 1649977179
transform 1 0 107916 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1173
timestamp 1649977179
transform 1 0 109020 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1185
timestamp 1649977179
transform 1 0 110124 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1197
timestamp 1649977179
transform 1 0 111228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1203
timestamp 1649977179
transform 1 0 111780 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1205
timestamp 1649977179
transform 1 0 111964 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1217
timestamp 1649977179
transform 1 0 113068 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1229
timestamp 1649977179
transform 1 0 114172 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1241
timestamp 1649977179
transform 1 0 115276 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1253
timestamp 1649977179
transform 1 0 116380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1259
timestamp 1649977179
transform 1 0 116932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_1261
timestamp 1649977179
transform 1 0 117116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_1273
timestamp 1649977179
transform 1 0 118220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_6
timestamp 1649977179
transform 1 0 1656 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_10
timestamp 1649977179
transform 1 0 2024 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_22
timestamp 1649977179
transform 1 0 3128 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_34
timestamp 1649977179
transform 1 0 4232 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_46
timestamp 1649977179
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1649977179
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1649977179
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1649977179
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1649977179
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1649977179
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1649977179
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1649977179
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1649977179
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1649977179
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1649977179
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1649977179
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1649977179
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1649977179
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_729
timestamp 1649977179
transform 1 0 68172 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_741
timestamp 1649977179
transform 1 0 69276 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_753
timestamp 1649977179
transform 1 0 70380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_765
timestamp 1649977179
transform 1 0 71484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 1649977179
transform 1 0 72588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 1649977179
transform 1 0 73140 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_785
timestamp 1649977179
transform 1 0 73324 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_797
timestamp 1649977179
transform 1 0 74428 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_809
timestamp 1649977179
transform 1 0 75532 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_821
timestamp 1649977179
transform 1 0 76636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_833
timestamp 1649977179
transform 1 0 77740 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_839
timestamp 1649977179
transform 1 0 78292 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_841
timestamp 1649977179
transform 1 0 78476 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_853
timestamp 1649977179
transform 1 0 79580 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_865
timestamp 1649977179
transform 1 0 80684 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_877
timestamp 1649977179
transform 1 0 81788 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_885
timestamp 1649977179
transform 1 0 82524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_890
timestamp 1649977179
transform 1 0 82984 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_897
timestamp 1649977179
transform 1 0 83628 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_909
timestamp 1649977179
transform 1 0 84732 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_921
timestamp 1649977179
transform 1 0 85836 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_933
timestamp 1649977179
transform 1 0 86940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_945
timestamp 1649977179
transform 1 0 88044 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_951
timestamp 1649977179
transform 1 0 88596 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_953
timestamp 1649977179
transform 1 0 88780 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_965
timestamp 1649977179
transform 1 0 89884 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_977
timestamp 1649977179
transform 1 0 90988 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_989
timestamp 1649977179
transform 1 0 92092 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1001
timestamp 1649977179
transform 1 0 93196 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1007
timestamp 1649977179
transform 1 0 93748 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1009
timestamp 1649977179
transform 1 0 93932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1021
timestamp 1649977179
transform 1 0 95036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1033
timestamp 1649977179
transform 1 0 96140 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1045
timestamp 1649977179
transform 1 0 97244 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1057
timestamp 1649977179
transform 1 0 98348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1063
timestamp 1649977179
transform 1 0 98900 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1065
timestamp 1649977179
transform 1 0 99084 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1077
timestamp 1649977179
transform 1 0 100188 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1089
timestamp 1649977179
transform 1 0 101292 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1101
timestamp 1649977179
transform 1 0 102396 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1113
timestamp 1649977179
transform 1 0 103500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1119
timestamp 1649977179
transform 1 0 104052 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1121
timestamp 1649977179
transform 1 0 104236 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1133
timestamp 1649977179
transform 1 0 105340 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1145
timestamp 1649977179
transform 1 0 106444 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1157
timestamp 1649977179
transform 1 0 107548 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1169
timestamp 1649977179
transform 1 0 108652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1175
timestamp 1649977179
transform 1 0 109204 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1177
timestamp 1649977179
transform 1 0 109388 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1189
timestamp 1649977179
transform 1 0 110492 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1201
timestamp 1649977179
transform 1 0 111596 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1213
timestamp 1649977179
transform 1 0 112700 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1225
timestamp 1649977179
transform 1 0 113804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1231
timestamp 1649977179
transform 1 0 114356 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1233
timestamp 1649977179
transform 1 0 114540 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1245
timestamp 1649977179
transform 1 0 115644 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1257
timestamp 1649977179
transform 1 0 116748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1269
timestamp 1649977179
transform 1 0 117852 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_349
timestamp 1649977179
transform 1 0 33212 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_359
timestamp 1649977179
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1649977179
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1649977179
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1649977179
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1649977179
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1649977179
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1649977179
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1649977179
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1649977179
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1649977179
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1649977179
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1649977179
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1649977179
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_725
timestamp 1649977179
transform 1 0 67804 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_737
timestamp 1649977179
transform 1 0 68908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 1649977179
transform 1 0 70012 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 1649977179
transform 1 0 70564 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_757
timestamp 1649977179
transform 1 0 70748 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_769
timestamp 1649977179
transform 1 0 71852 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_781
timestamp 1649977179
transform 1 0 72956 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_793
timestamp 1649977179
transform 1 0 74060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 1649977179
transform 1 0 75164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 1649977179
transform 1 0 75716 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_813
timestamp 1649977179
transform 1 0 75900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_825
timestamp 1649977179
transform 1 0 77004 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_837
timestamp 1649977179
transform 1 0 78108 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_849
timestamp 1649977179
transform 1 0 79212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_861
timestamp 1649977179
transform 1 0 80316 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_867
timestamp 1649977179
transform 1 0 80868 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_869
timestamp 1649977179
transform 1 0 81052 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_881
timestamp 1649977179
transform 1 0 82156 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_893
timestamp 1649977179
transform 1 0 83260 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_905
timestamp 1649977179
transform 1 0 84364 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_917
timestamp 1649977179
transform 1 0 85468 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_923
timestamp 1649977179
transform 1 0 86020 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_925
timestamp 1649977179
transform 1 0 86204 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_937
timestamp 1649977179
transform 1 0 87308 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_949
timestamp 1649977179
transform 1 0 88412 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_961
timestamp 1649977179
transform 1 0 89516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_973
timestamp 1649977179
transform 1 0 90620 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_979
timestamp 1649977179
transform 1 0 91172 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_981
timestamp 1649977179
transform 1 0 91356 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_993
timestamp 1649977179
transform 1 0 92460 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1005
timestamp 1649977179
transform 1 0 93564 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1017
timestamp 1649977179
transform 1 0 94668 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1029
timestamp 1649977179
transform 1 0 95772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1035
timestamp 1649977179
transform 1 0 96324 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1037
timestamp 1649977179
transform 1 0 96508 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1049
timestamp 1649977179
transform 1 0 97612 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1061
timestamp 1649977179
transform 1 0 98716 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1073
timestamp 1649977179
transform 1 0 99820 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1085
timestamp 1649977179
transform 1 0 100924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1091
timestamp 1649977179
transform 1 0 101476 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1093
timestamp 1649977179
transform 1 0 101660 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1105
timestamp 1649977179
transform 1 0 102764 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1117
timestamp 1649977179
transform 1 0 103868 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1129
timestamp 1649977179
transform 1 0 104972 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1141
timestamp 1649977179
transform 1 0 106076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1147
timestamp 1649977179
transform 1 0 106628 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1149
timestamp 1649977179
transform 1 0 106812 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1161
timestamp 1649977179
transform 1 0 107916 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1173
timestamp 1649977179
transform 1 0 109020 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1185
timestamp 1649977179
transform 1 0 110124 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1197
timestamp 1649977179
transform 1 0 111228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1203
timestamp 1649977179
transform 1 0 111780 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1205
timestamp 1649977179
transform 1 0 111964 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1217
timestamp 1649977179
transform 1 0 113068 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1229
timestamp 1649977179
transform 1 0 114172 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1241
timestamp 1649977179
transform 1 0 115276 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1253
timestamp 1649977179
transform 1 0 116380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1259
timestamp 1649977179
transform 1 0 116932 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1261
timestamp 1649977179
transform 1 0 117116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_1273
timestamp 1649977179
transform 1 0 118220 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_345
timestamp 1649977179
transform 1 0 32844 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_357
timestamp 1649977179
transform 1 0 33948 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_369
timestamp 1649977179
transform 1 0 35052 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_381
timestamp 1649977179
transform 1 0 36156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1649977179
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1649977179
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1649977179
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1649977179
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1649977179
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1649977179
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1649977179
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1649977179
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1649977179
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1649977179
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1649977179
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1649977179
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_729
timestamp 1649977179
transform 1 0 68172 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_741
timestamp 1649977179
transform 1 0 69276 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_753
timestamp 1649977179
transform 1 0 70380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_765
timestamp 1649977179
transform 1 0 71484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 1649977179
transform 1 0 72588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 1649977179
transform 1 0 73140 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_785
timestamp 1649977179
transform 1 0 73324 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_797
timestamp 1649977179
transform 1 0 74428 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_809
timestamp 1649977179
transform 1 0 75532 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_821
timestamp 1649977179
transform 1 0 76636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_833
timestamp 1649977179
transform 1 0 77740 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_839
timestamp 1649977179
transform 1 0 78292 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_841
timestamp 1649977179
transform 1 0 78476 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_853
timestamp 1649977179
transform 1 0 79580 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_865
timestamp 1649977179
transform 1 0 80684 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_877
timestamp 1649977179
transform 1 0 81788 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_889
timestamp 1649977179
transform 1 0 82892 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_895
timestamp 1649977179
transform 1 0 83444 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_897
timestamp 1649977179
transform 1 0 83628 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_909
timestamp 1649977179
transform 1 0 84732 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_921
timestamp 1649977179
transform 1 0 85836 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_933
timestamp 1649977179
transform 1 0 86940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_945
timestamp 1649977179
transform 1 0 88044 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_951
timestamp 1649977179
transform 1 0 88596 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_953
timestamp 1649977179
transform 1 0 88780 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_965
timestamp 1649977179
transform 1 0 89884 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_977
timestamp 1649977179
transform 1 0 90988 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_989
timestamp 1649977179
transform 1 0 92092 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1001
timestamp 1649977179
transform 1 0 93196 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1007
timestamp 1649977179
transform 1 0 93748 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1009
timestamp 1649977179
transform 1 0 93932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1021
timestamp 1649977179
transform 1 0 95036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1033
timestamp 1649977179
transform 1 0 96140 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1045
timestamp 1649977179
transform 1 0 97244 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1057
timestamp 1649977179
transform 1 0 98348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1063
timestamp 1649977179
transform 1 0 98900 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1065
timestamp 1649977179
transform 1 0 99084 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1077
timestamp 1649977179
transform 1 0 100188 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1089
timestamp 1649977179
transform 1 0 101292 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1101
timestamp 1649977179
transform 1 0 102396 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1113
timestamp 1649977179
transform 1 0 103500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1119
timestamp 1649977179
transform 1 0 104052 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1121
timestamp 1649977179
transform 1 0 104236 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1133
timestamp 1649977179
transform 1 0 105340 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1145
timestamp 1649977179
transform 1 0 106444 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1157
timestamp 1649977179
transform 1 0 107548 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1169
timestamp 1649977179
transform 1 0 108652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1175
timestamp 1649977179
transform 1 0 109204 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1177
timestamp 1649977179
transform 1 0 109388 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1189
timestamp 1649977179
transform 1 0 110492 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1201
timestamp 1649977179
transform 1 0 111596 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1213
timestamp 1649977179
transform 1 0 112700 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1225
timestamp 1649977179
transform 1 0 113804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1231
timestamp 1649977179
transform 1 0 114356 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1233
timestamp 1649977179
transform 1 0 114540 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1245
timestamp 1649977179
transform 1 0 115644 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1257
timestamp 1649977179
transform 1 0 116748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_1273
timestamp 1649977179
transform 1 0 118220 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_6
timestamp 1649977179
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_18
timestamp 1649977179
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1649977179
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1649977179
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1649977179
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1649977179
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1649977179
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1649977179
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1649977179
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1649977179
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1649977179
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1649977179
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1649977179
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1649977179
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_725
timestamp 1649977179
transform 1 0 67804 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_737
timestamp 1649977179
transform 1 0 68908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 1649977179
transform 1 0 70012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 1649977179
transform 1 0 70564 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_757
timestamp 1649977179
transform 1 0 70748 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_769
timestamp 1649977179
transform 1 0 71852 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_781
timestamp 1649977179
transform 1 0 72956 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_793
timestamp 1649977179
transform 1 0 74060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 1649977179
transform 1 0 75164 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 1649977179
transform 1 0 75716 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_813
timestamp 1649977179
transform 1 0 75900 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_825
timestamp 1649977179
transform 1 0 77004 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_837
timestamp 1649977179
transform 1 0 78108 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_849
timestamp 1649977179
transform 1 0 79212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_861
timestamp 1649977179
transform 1 0 80316 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_867
timestamp 1649977179
transform 1 0 80868 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_869
timestamp 1649977179
transform 1 0 81052 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_881
timestamp 1649977179
transform 1 0 82156 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_893
timestamp 1649977179
transform 1 0 83260 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_905
timestamp 1649977179
transform 1 0 84364 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_917
timestamp 1649977179
transform 1 0 85468 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_923
timestamp 1649977179
transform 1 0 86020 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_925
timestamp 1649977179
transform 1 0 86204 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_937
timestamp 1649977179
transform 1 0 87308 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_949
timestamp 1649977179
transform 1 0 88412 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_961
timestamp 1649977179
transform 1 0 89516 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_973
timestamp 1649977179
transform 1 0 90620 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_979
timestamp 1649977179
transform 1 0 91172 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_981
timestamp 1649977179
transform 1 0 91356 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_993
timestamp 1649977179
transform 1 0 92460 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1005
timestamp 1649977179
transform 1 0 93564 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1017
timestamp 1649977179
transform 1 0 94668 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1029
timestamp 1649977179
transform 1 0 95772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1035
timestamp 1649977179
transform 1 0 96324 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1037
timestamp 1649977179
transform 1 0 96508 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1049
timestamp 1649977179
transform 1 0 97612 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1061
timestamp 1649977179
transform 1 0 98716 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1073
timestamp 1649977179
transform 1 0 99820 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1085
timestamp 1649977179
transform 1 0 100924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1091
timestamp 1649977179
transform 1 0 101476 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1093
timestamp 1649977179
transform 1 0 101660 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1105
timestamp 1649977179
transform 1 0 102764 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1117
timestamp 1649977179
transform 1 0 103868 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1129
timestamp 1649977179
transform 1 0 104972 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1141
timestamp 1649977179
transform 1 0 106076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1147
timestamp 1649977179
transform 1 0 106628 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1149
timestamp 1649977179
transform 1 0 106812 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1161
timestamp 1649977179
transform 1 0 107916 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1173
timestamp 1649977179
transform 1 0 109020 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1185
timestamp 1649977179
transform 1 0 110124 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1197
timestamp 1649977179
transform 1 0 111228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1203
timestamp 1649977179
transform 1 0 111780 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1205
timestamp 1649977179
transform 1 0 111964 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1217
timestamp 1649977179
transform 1 0 113068 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1229
timestamp 1649977179
transform 1 0 114172 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1241
timestamp 1649977179
transform 1 0 115276 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1253
timestamp 1649977179
transform 1 0 116380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1259
timestamp 1649977179
transform 1 0 116932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_1261
timestamp 1649977179
transform 1 0 117116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_1273
timestamp 1649977179
transform 1 0 118220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_25
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_37
timestamp 1649977179
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1649977179
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1649977179
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1649977179
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1649977179
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1649977179
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1649977179
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1649977179
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1649977179
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1649977179
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1649977179
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1649977179
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1649977179
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_729
timestamp 1649977179
transform 1 0 68172 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_741
timestamp 1649977179
transform 1 0 69276 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_753
timestamp 1649977179
transform 1 0 70380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_765
timestamp 1649977179
transform 1 0 71484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 1649977179
transform 1 0 72588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 1649977179
transform 1 0 73140 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_785
timestamp 1649977179
transform 1 0 73324 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_797
timestamp 1649977179
transform 1 0 74428 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_809
timestamp 1649977179
transform 1 0 75532 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_821
timestamp 1649977179
transform 1 0 76636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_833
timestamp 1649977179
transform 1 0 77740 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_839
timestamp 1649977179
transform 1 0 78292 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_841
timestamp 1649977179
transform 1 0 78476 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_853
timestamp 1649977179
transform 1 0 79580 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_865
timestamp 1649977179
transform 1 0 80684 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_877
timestamp 1649977179
transform 1 0 81788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_889
timestamp 1649977179
transform 1 0 82892 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_895
timestamp 1649977179
transform 1 0 83444 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_897
timestamp 1649977179
transform 1 0 83628 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_909
timestamp 1649977179
transform 1 0 84732 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_921
timestamp 1649977179
transform 1 0 85836 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_933
timestamp 1649977179
transform 1 0 86940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_945
timestamp 1649977179
transform 1 0 88044 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_951
timestamp 1649977179
transform 1 0 88596 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_953
timestamp 1649977179
transform 1 0 88780 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_965
timestamp 1649977179
transform 1 0 89884 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_977
timestamp 1649977179
transform 1 0 90988 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_989
timestamp 1649977179
transform 1 0 92092 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1001
timestamp 1649977179
transform 1 0 93196 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1007
timestamp 1649977179
transform 1 0 93748 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1009
timestamp 1649977179
transform 1 0 93932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1021
timestamp 1649977179
transform 1 0 95036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1033
timestamp 1649977179
transform 1 0 96140 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1045
timestamp 1649977179
transform 1 0 97244 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1057
timestamp 1649977179
transform 1 0 98348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1063
timestamp 1649977179
transform 1 0 98900 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1065
timestamp 1649977179
transform 1 0 99084 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1077
timestamp 1649977179
transform 1 0 100188 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1089
timestamp 1649977179
transform 1 0 101292 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1101
timestamp 1649977179
transform 1 0 102396 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1113
timestamp 1649977179
transform 1 0 103500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1119
timestamp 1649977179
transform 1 0 104052 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1121
timestamp 1649977179
transform 1 0 104236 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1133
timestamp 1649977179
transform 1 0 105340 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1145
timestamp 1649977179
transform 1 0 106444 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1157
timestamp 1649977179
transform 1 0 107548 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1169
timestamp 1649977179
transform 1 0 108652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1175
timestamp 1649977179
transform 1 0 109204 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1177
timestamp 1649977179
transform 1 0 109388 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1189
timestamp 1649977179
transform 1 0 110492 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1201
timestamp 1649977179
transform 1 0 111596 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1213
timestamp 1649977179
transform 1 0 112700 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1225
timestamp 1649977179
transform 1 0 113804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1231
timestamp 1649977179
transform 1 0 114356 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1233
timestamp 1649977179
transform 1 0 114540 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1245
timestamp 1649977179
transform 1 0 115644 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1257
timestamp 1649977179
transform 1 0 116748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_1269
timestamp 1649977179
transform 1 0 117852 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_6
timestamp 1649977179
transform 1 0 1656 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp 1649977179
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1649977179
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1649977179
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1649977179
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1649977179
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1649977179
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1649977179
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1649977179
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1649977179
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1649977179
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1649977179
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1649977179
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_725
timestamp 1649977179
transform 1 0 67804 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_737
timestamp 1649977179
transform 1 0 68908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 1649977179
transform 1 0 70012 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 1649977179
transform 1 0 70564 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_757
timestamp 1649977179
transform 1 0 70748 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_769
timestamp 1649977179
transform 1 0 71852 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_781
timestamp 1649977179
transform 1 0 72956 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_793
timestamp 1649977179
transform 1 0 74060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 1649977179
transform 1 0 75164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 1649977179
transform 1 0 75716 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_813
timestamp 1649977179
transform 1 0 75900 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_825
timestamp 1649977179
transform 1 0 77004 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_837
timestamp 1649977179
transform 1 0 78108 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_853
timestamp 1649977179
transform 1 0 79580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_860
timestamp 1649977179
transform 1 0 80224 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_869
timestamp 1649977179
transform 1 0 81052 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_881
timestamp 1649977179
transform 1 0 82156 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_893
timestamp 1649977179
transform 1 0 83260 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_905
timestamp 1649977179
transform 1 0 84364 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_917
timestamp 1649977179
transform 1 0 85468 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_923
timestamp 1649977179
transform 1 0 86020 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_925
timestamp 1649977179
transform 1 0 86204 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_937
timestamp 1649977179
transform 1 0 87308 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_949
timestamp 1649977179
transform 1 0 88412 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_961
timestamp 1649977179
transform 1 0 89516 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_973
timestamp 1649977179
transform 1 0 90620 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_979
timestamp 1649977179
transform 1 0 91172 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_981
timestamp 1649977179
transform 1 0 91356 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_993
timestamp 1649977179
transform 1 0 92460 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1005
timestamp 1649977179
transform 1 0 93564 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1017
timestamp 1649977179
transform 1 0 94668 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1029
timestamp 1649977179
transform 1 0 95772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1035
timestamp 1649977179
transform 1 0 96324 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1037
timestamp 1649977179
transform 1 0 96508 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1049
timestamp 1649977179
transform 1 0 97612 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1061
timestamp 1649977179
transform 1 0 98716 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1073
timestamp 1649977179
transform 1 0 99820 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1085
timestamp 1649977179
transform 1 0 100924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1091
timestamp 1649977179
transform 1 0 101476 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1093
timestamp 1649977179
transform 1 0 101660 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1105
timestamp 1649977179
transform 1 0 102764 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1117
timestamp 1649977179
transform 1 0 103868 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1129
timestamp 1649977179
transform 1 0 104972 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1141
timestamp 1649977179
transform 1 0 106076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1147
timestamp 1649977179
transform 1 0 106628 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1149
timestamp 1649977179
transform 1 0 106812 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1161
timestamp 1649977179
transform 1 0 107916 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1173
timestamp 1649977179
transform 1 0 109020 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1185
timestamp 1649977179
transform 1 0 110124 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1197
timestamp 1649977179
transform 1 0 111228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1203
timestamp 1649977179
transform 1 0 111780 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1205
timestamp 1649977179
transform 1 0 111964 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_1217
timestamp 1649977179
transform 1 0 113068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1221
timestamp 1649977179
transform 1 0 113436 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1226
timestamp 1649977179
transform 1 0 113896 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1238
timestamp 1649977179
transform 1 0 115000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_1250
timestamp 1649977179
transform 1 0 116104 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_1258
timestamp 1649977179
transform 1 0 116840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_1261
timestamp 1649977179
transform 1 0 117116 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1269
timestamp 1649977179
transform 1 0 117852 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_1273
timestamp 1649977179
transform 1 0 118220 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1649977179
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1649977179
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1649977179
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1649977179
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1649977179
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1649977179
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1649977179
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1649977179
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1649977179
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1649977179
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1649977179
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_729
timestamp 1649977179
transform 1 0 68172 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_741
timestamp 1649977179
transform 1 0 69276 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_753
timestamp 1649977179
transform 1 0 70380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_765
timestamp 1649977179
transform 1 0 71484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_773
timestamp 1649977179
transform 1 0 72220 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_781
timestamp 1649977179
transform 1 0 72956 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_785
timestamp 1649977179
transform 1 0 73324 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_797
timestamp 1649977179
transform 1 0 74428 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_809
timestamp 1649977179
transform 1 0 75532 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_821
timestamp 1649977179
transform 1 0 76636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_833
timestamp 1649977179
transform 1 0 77740 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_839
timestamp 1649977179
transform 1 0 78292 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_841
timestamp 1649977179
transform 1 0 78476 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_852
timestamp 1649977179
transform 1 0 79488 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_856
timestamp 1649977179
transform 1 0 79856 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_868
timestamp 1649977179
transform 1 0 80960 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_880
timestamp 1649977179
transform 1 0 82064 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_892
timestamp 1649977179
transform 1 0 83168 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_907
timestamp 1649977179
transform 1 0 84548 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_919
timestamp 1649977179
transform 1 0 85652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_931
timestamp 1649977179
transform 1 0 86756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_943
timestamp 1649977179
transform 1 0 87860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_951
timestamp 1649977179
transform 1 0 88596 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_953
timestamp 1649977179
transform 1 0 88780 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_965
timestamp 1649977179
transform 1 0 89884 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_977
timestamp 1649977179
transform 1 0 90988 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_989
timestamp 1649977179
transform 1 0 92092 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1001
timestamp 1649977179
transform 1 0 93196 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1007
timestamp 1649977179
transform 1 0 93748 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1009
timestamp 1649977179
transform 1 0 93932 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1021
timestamp 1649977179
transform 1 0 95036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1033
timestamp 1649977179
transform 1 0 96140 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1045
timestamp 1649977179
transform 1 0 97244 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1057
timestamp 1649977179
transform 1 0 98348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1063
timestamp 1649977179
transform 1 0 98900 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1065
timestamp 1649977179
transform 1 0 99084 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1077
timestamp 1649977179
transform 1 0 100188 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1089
timestamp 1649977179
transform 1 0 101292 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1101
timestamp 1649977179
transform 1 0 102396 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1113
timestamp 1649977179
transform 1 0 103500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1119
timestamp 1649977179
transform 1 0 104052 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1121
timestamp 1649977179
transform 1 0 104236 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1133
timestamp 1649977179
transform 1 0 105340 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1145
timestamp 1649977179
transform 1 0 106444 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1157
timestamp 1649977179
transform 1 0 107548 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1169
timestamp 1649977179
transform 1 0 108652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1175
timestamp 1649977179
transform 1 0 109204 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1177
timestamp 1649977179
transform 1 0 109388 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1189
timestamp 1649977179
transform 1 0 110492 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1201
timestamp 1649977179
transform 1 0 111596 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1213
timestamp 1649977179
transform 1 0 112700 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1225
timestamp 1649977179
transform 1 0 113804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1231
timestamp 1649977179
transform 1 0 114356 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1236
timestamp 1649977179
transform 1 0 114816 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1248
timestamp 1649977179
transform 1 0 115920 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1260
timestamp 1649977179
transform 1 0 117024 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_1272
timestamp 1649977179
transform 1 0 118128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1276
timestamp 1649977179
transform 1 0 118496 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_577
timestamp 1649977179
transform 1 0 54188 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_584
timestamp 1649977179
transform 1 0 54832 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_599
timestamp 1649977179
transform 1 0 56212 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_611
timestamp 1649977179
transform 1 0 57316 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_623
timestamp 1649977179
transform 1 0 58420 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_635
timestamp 1649977179
transform 1 0 59524 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1649977179
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1649977179
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1649977179
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1649977179
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1649977179
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1649977179
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1649977179
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1649977179
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1649977179
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_725
timestamp 1649977179
transform 1 0 67804 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_737
timestamp 1649977179
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 1649977179
transform 1 0 70012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 1649977179
transform 1 0 70564 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_757
timestamp 1649977179
transform 1 0 70748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_769
timestamp 1649977179
transform 1 0 71852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_773
timestamp 1649977179
transform 1 0 72220 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_783
timestamp 1649977179
transform 1 0 73140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_795
timestamp 1649977179
transform 1 0 74244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_807
timestamp 1649977179
transform 1 0 75348 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 1649977179
transform 1 0 75716 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_813
timestamp 1649977179
transform 1 0 75900 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_825
timestamp 1649977179
transform 1 0 77004 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_837
timestamp 1649977179
transform 1 0 78108 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_849
timestamp 1649977179
transform 1 0 79212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_861
timestamp 1649977179
transform 1 0 80316 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_867
timestamp 1649977179
transform 1 0 80868 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_869
timestamp 1649977179
transform 1 0 81052 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_881
timestamp 1649977179
transform 1 0 82156 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_893
timestamp 1649977179
transform 1 0 83260 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_901
timestamp 1649977179
transform 1 0 83996 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_904
timestamp 1649977179
transform 1 0 84272 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_915
timestamp 1649977179
transform 1 0 85284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_923
timestamp 1649977179
transform 1 0 86020 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_925
timestamp 1649977179
transform 1 0 86204 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_937
timestamp 1649977179
transform 1 0 87308 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_949
timestamp 1649977179
transform 1 0 88412 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_961
timestamp 1649977179
transform 1 0 89516 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_973
timestamp 1649977179
transform 1 0 90620 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_979
timestamp 1649977179
transform 1 0 91172 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_981
timestamp 1649977179
transform 1 0 91356 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_993
timestamp 1649977179
transform 1 0 92460 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1005
timestamp 1649977179
transform 1 0 93564 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1017
timestamp 1649977179
transform 1 0 94668 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1029
timestamp 1649977179
transform 1 0 95772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1035
timestamp 1649977179
transform 1 0 96324 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1037
timestamp 1649977179
transform 1 0 96508 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1049
timestamp 1649977179
transform 1 0 97612 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1061
timestamp 1649977179
transform 1 0 98716 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1073
timestamp 1649977179
transform 1 0 99820 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1085
timestamp 1649977179
transform 1 0 100924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1091
timestamp 1649977179
transform 1 0 101476 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1093
timestamp 1649977179
transform 1 0 101660 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1105
timestamp 1649977179
transform 1 0 102764 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1117
timestamp 1649977179
transform 1 0 103868 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1129
timestamp 1649977179
transform 1 0 104972 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1141
timestamp 1649977179
transform 1 0 106076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1147
timestamp 1649977179
transform 1 0 106628 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1149
timestamp 1649977179
transform 1 0 106812 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1161
timestamp 1649977179
transform 1 0 107916 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1173
timestamp 1649977179
transform 1 0 109020 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1185
timestamp 1649977179
transform 1 0 110124 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1197
timestamp 1649977179
transform 1 0 111228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1203
timestamp 1649977179
transform 1 0 111780 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1205
timestamp 1649977179
transform 1 0 111964 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1217
timestamp 1649977179
transform 1 0 113068 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1229
timestamp 1649977179
transform 1 0 114172 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1241
timestamp 1649977179
transform 1 0 115276 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1253
timestamp 1649977179
transform 1 0 116380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1259
timestamp 1649977179
transform 1 0 116932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_1261
timestamp 1649977179
transform 1 0 117116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1269
timestamp 1649977179
transform 1 0 117852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_1273
timestamp 1649977179
transform 1 0 118220 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_7
timestamp 1649977179
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_19
timestamp 1649977179
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_31
timestamp 1649977179
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1649977179
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_509
timestamp 1649977179
transform 1 0 47932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_521
timestamp 1649977179
transform 1 0 49036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_533
timestamp 1649977179
transform 1 0 50140 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_545
timestamp 1649977179
transform 1 0 51244 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_557
timestamp 1649977179
transform 1 0 52348 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1649977179
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1649977179
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1649977179
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1649977179
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1649977179
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1649977179
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1649977179
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1649977179
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1649977179
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1649977179
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1649977179
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_738
timestamp 1649977179
transform 1 0 69000 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_750
timestamp 1649977179
transform 1 0 70104 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_762
timestamp 1649977179
transform 1 0 71208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_774
timestamp 1649977179
transform 1 0 72312 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_782
timestamp 1649977179
transform 1 0 73048 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_785
timestamp 1649977179
transform 1 0 73324 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_797
timestamp 1649977179
transform 1 0 74428 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_809
timestamp 1649977179
transform 1 0 75532 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_821
timestamp 1649977179
transform 1 0 76636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_833
timestamp 1649977179
transform 1 0 77740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_839
timestamp 1649977179
transform 1 0 78292 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_841
timestamp 1649977179
transform 1 0 78476 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_853
timestamp 1649977179
transform 1 0 79580 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_865
timestamp 1649977179
transform 1 0 80684 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_877
timestamp 1649977179
transform 1 0 81788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_889
timestamp 1649977179
transform 1 0 82892 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_895
timestamp 1649977179
transform 1 0 83444 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_897
timestamp 1649977179
transform 1 0 83628 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_909
timestamp 1649977179
transform 1 0 84732 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_921
timestamp 1649977179
transform 1 0 85836 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_933
timestamp 1649977179
transform 1 0 86940 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_945
timestamp 1649977179
transform 1 0 88044 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_951
timestamp 1649977179
transform 1 0 88596 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_953
timestamp 1649977179
transform 1 0 88780 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_965
timestamp 1649977179
transform 1 0 89884 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_977
timestamp 1649977179
transform 1 0 90988 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_989
timestamp 1649977179
transform 1 0 92092 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1001
timestamp 1649977179
transform 1 0 93196 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1007
timestamp 1649977179
transform 1 0 93748 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1009
timestamp 1649977179
transform 1 0 93932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1021
timestamp 1649977179
transform 1 0 95036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1033
timestamp 1649977179
transform 1 0 96140 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1045
timestamp 1649977179
transform 1 0 97244 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1057
timestamp 1649977179
transform 1 0 98348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1063
timestamp 1649977179
transform 1 0 98900 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1065
timestamp 1649977179
transform 1 0 99084 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1077
timestamp 1649977179
transform 1 0 100188 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1089
timestamp 1649977179
transform 1 0 101292 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1101
timestamp 1649977179
transform 1 0 102396 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1113
timestamp 1649977179
transform 1 0 103500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1119
timestamp 1649977179
transform 1 0 104052 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1121
timestamp 1649977179
transform 1 0 104236 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1133
timestamp 1649977179
transform 1 0 105340 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1145
timestamp 1649977179
transform 1 0 106444 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1157
timestamp 1649977179
transform 1 0 107548 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1169
timestamp 1649977179
transform 1 0 108652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1175
timestamp 1649977179
transform 1 0 109204 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1177
timestamp 1649977179
transform 1 0 109388 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1189
timestamp 1649977179
transform 1 0 110492 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1201
timestamp 1649977179
transform 1 0 111596 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1213
timestamp 1649977179
transform 1 0 112700 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1225
timestamp 1649977179
transform 1 0 113804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1231
timestamp 1649977179
transform 1 0 114356 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1233
timestamp 1649977179
transform 1 0 114540 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1245
timestamp 1649977179
transform 1 0 115644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1257
timestamp 1649977179
transform 1 0 116748 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_1273
timestamp 1649977179
transform 1 0 118220 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_6
timestamp 1649977179
transform 1 0 1656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_18
timestamp 1649977179
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1649977179
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1649977179
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_521
timestamp 1649977179
transform 1 0 49036 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_527
timestamp 1649977179
transform 1 0 49588 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_542
timestamp 1649977179
transform 1 0 50968 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_554
timestamp 1649977179
transform 1 0 52072 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_566
timestamp 1649977179
transform 1 0 53176 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_578
timestamp 1649977179
transform 1 0 54280 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_586
timestamp 1649977179
transform 1 0 55016 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1649977179
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1649977179
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1649977179
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1649977179
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1649977179
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1649977179
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1649977179
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1649977179
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1649977179
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1649977179
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1649977179
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_725
timestamp 1649977179
transform 1 0 67804 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_731
timestamp 1649977179
transform 1 0 68356 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_736
timestamp 1649977179
transform 1 0 68816 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_748
timestamp 1649977179
transform 1 0 69920 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_757
timestamp 1649977179
transform 1 0 70748 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_769
timestamp 1649977179
transform 1 0 71852 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_781
timestamp 1649977179
transform 1 0 72956 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_793
timestamp 1649977179
transform 1 0 74060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 1649977179
transform 1 0 75164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 1649977179
transform 1 0 75716 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_813
timestamp 1649977179
transform 1 0 75900 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_825
timestamp 1649977179
transform 1 0 77004 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_837
timestamp 1649977179
transform 1 0 78108 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_849
timestamp 1649977179
transform 1 0 79212 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_861
timestamp 1649977179
transform 1 0 80316 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_867
timestamp 1649977179
transform 1 0 80868 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_869
timestamp 1649977179
transform 1 0 81052 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_881
timestamp 1649977179
transform 1 0 82156 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_893
timestamp 1649977179
transform 1 0 83260 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_905
timestamp 1649977179
transform 1 0 84364 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_917
timestamp 1649977179
transform 1 0 85468 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_923
timestamp 1649977179
transform 1 0 86020 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_925
timestamp 1649977179
transform 1 0 86204 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_937
timestamp 1649977179
transform 1 0 87308 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_949
timestamp 1649977179
transform 1 0 88412 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_961
timestamp 1649977179
transform 1 0 89516 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_973
timestamp 1649977179
transform 1 0 90620 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_979
timestamp 1649977179
transform 1 0 91172 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_981
timestamp 1649977179
transform 1 0 91356 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_993
timestamp 1649977179
transform 1 0 92460 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1005
timestamp 1649977179
transform 1 0 93564 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1017
timestamp 1649977179
transform 1 0 94668 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1029
timestamp 1649977179
transform 1 0 95772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1035
timestamp 1649977179
transform 1 0 96324 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1037
timestamp 1649977179
transform 1 0 96508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1049
timestamp 1649977179
transform 1 0 97612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1061
timestamp 1649977179
transform 1 0 98716 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1073
timestamp 1649977179
transform 1 0 99820 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1085
timestamp 1649977179
transform 1 0 100924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1091
timestamp 1649977179
transform 1 0 101476 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1093
timestamp 1649977179
transform 1 0 101660 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1105
timestamp 1649977179
transform 1 0 102764 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1117
timestamp 1649977179
transform 1 0 103868 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1129
timestamp 1649977179
transform 1 0 104972 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1141
timestamp 1649977179
transform 1 0 106076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1147
timestamp 1649977179
transform 1 0 106628 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1149
timestamp 1649977179
transform 1 0 106812 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1161
timestamp 1649977179
transform 1 0 107916 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1173
timestamp 1649977179
transform 1 0 109020 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1185
timestamp 1649977179
transform 1 0 110124 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1197
timestamp 1649977179
transform 1 0 111228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1203
timestamp 1649977179
transform 1 0 111780 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1205
timestamp 1649977179
transform 1 0 111964 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1217
timestamp 1649977179
transform 1 0 113068 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1229
timestamp 1649977179
transform 1 0 114172 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1241
timestamp 1649977179
transform 1 0 115276 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1253
timestamp 1649977179
transform 1 0 116380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1259
timestamp 1649977179
transform 1 0 116932 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1261
timestamp 1649977179
transform 1 0 117116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_1273
timestamp 1649977179
transform 1 0 118220 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1649977179
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1649977179
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1649977179
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1649977179
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1649977179
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1649977179
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1649977179
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1649977179
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1649977179
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1649977179
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1649977179
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_729
timestamp 1649977179
transform 1 0 68172 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_741
timestamp 1649977179
transform 1 0 69276 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_753
timestamp 1649977179
transform 1 0 70380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_765
timestamp 1649977179
transform 1 0 71484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 1649977179
transform 1 0 72588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 1649977179
transform 1 0 73140 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_785
timestamp 1649977179
transform 1 0 73324 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_797
timestamp 1649977179
transform 1 0 74428 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_809
timestamp 1649977179
transform 1 0 75532 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_821
timestamp 1649977179
transform 1 0 76636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_833
timestamp 1649977179
transform 1 0 77740 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_839
timestamp 1649977179
transform 1 0 78292 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_841
timestamp 1649977179
transform 1 0 78476 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_853
timestamp 1649977179
transform 1 0 79580 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_865
timestamp 1649977179
transform 1 0 80684 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_877
timestamp 1649977179
transform 1 0 81788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_889
timestamp 1649977179
transform 1 0 82892 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_895
timestamp 1649977179
transform 1 0 83444 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_897
timestamp 1649977179
transform 1 0 83628 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_909
timestamp 1649977179
transform 1 0 84732 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_921
timestamp 1649977179
transform 1 0 85836 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_933
timestamp 1649977179
transform 1 0 86940 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_945
timestamp 1649977179
transform 1 0 88044 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_951
timestamp 1649977179
transform 1 0 88596 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_953
timestamp 1649977179
transform 1 0 88780 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_965
timestamp 1649977179
transform 1 0 89884 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_977
timestamp 1649977179
transform 1 0 90988 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_989
timestamp 1649977179
transform 1 0 92092 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1001
timestamp 1649977179
transform 1 0 93196 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1007
timestamp 1649977179
transform 1 0 93748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_1009
timestamp 1649977179
transform 1 0 93932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1013
timestamp 1649977179
transform 1 0 94300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_1023
timestamp 1649977179
transform 1 0 95220 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1030
timestamp 1649977179
transform 1 0 95864 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1042
timestamp 1649977179
transform 1 0 96968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1054
timestamp 1649977179
transform 1 0 98072 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_1062
timestamp 1649977179
transform 1 0 98808 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1065
timestamp 1649977179
transform 1 0 99084 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1077
timestamp 1649977179
transform 1 0 100188 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1089
timestamp 1649977179
transform 1 0 101292 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1101
timestamp 1649977179
transform 1 0 102396 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1113
timestamp 1649977179
transform 1 0 103500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1119
timestamp 1649977179
transform 1 0 104052 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1121
timestamp 1649977179
transform 1 0 104236 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1133
timestamp 1649977179
transform 1 0 105340 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1145
timestamp 1649977179
transform 1 0 106444 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1157
timestamp 1649977179
transform 1 0 107548 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1169
timestamp 1649977179
transform 1 0 108652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1175
timestamp 1649977179
transform 1 0 109204 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1177
timestamp 1649977179
transform 1 0 109388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1189
timestamp 1649977179
transform 1 0 110492 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1201
timestamp 1649977179
transform 1 0 111596 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1213
timestamp 1649977179
transform 1 0 112700 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1225
timestamp 1649977179
transform 1 0 113804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1231
timestamp 1649977179
transform 1 0 114356 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1233
timestamp 1649977179
transform 1 0 114540 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1245
timestamp 1649977179
transform 1 0 115644 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1257
timestamp 1649977179
transform 1 0 116748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1269
timestamp 1649977179
transform 1 0 117852 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_1273
timestamp 1649977179
transform 1 0 118220 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1649977179
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1649977179
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1649977179
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1649977179
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1649977179
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1649977179
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1649977179
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1649977179
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1649977179
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1649977179
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1649977179
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_725
timestamp 1649977179
transform 1 0 67804 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_737
timestamp 1649977179
transform 1 0 68908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 1649977179
transform 1 0 70012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 1649977179
transform 1 0 70564 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_757
timestamp 1649977179
transform 1 0 70748 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_769
timestamp 1649977179
transform 1 0 71852 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_781
timestamp 1649977179
transform 1 0 72956 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_793
timestamp 1649977179
transform 1 0 74060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 1649977179
transform 1 0 75164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 1649977179
transform 1 0 75716 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_813
timestamp 1649977179
transform 1 0 75900 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_825
timestamp 1649977179
transform 1 0 77004 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_837
timestamp 1649977179
transform 1 0 78108 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_849
timestamp 1649977179
transform 1 0 79212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_861
timestamp 1649977179
transform 1 0 80316 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_867
timestamp 1649977179
transform 1 0 80868 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_869
timestamp 1649977179
transform 1 0 81052 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_881
timestamp 1649977179
transform 1 0 82156 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_893
timestamp 1649977179
transform 1 0 83260 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_905
timestamp 1649977179
transform 1 0 84364 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_917
timestamp 1649977179
transform 1 0 85468 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_923
timestamp 1649977179
transform 1 0 86020 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_925
timestamp 1649977179
transform 1 0 86204 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_937
timestamp 1649977179
transform 1 0 87308 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_949
timestamp 1649977179
transform 1 0 88412 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_961
timestamp 1649977179
transform 1 0 89516 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_973
timestamp 1649977179
transform 1 0 90620 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_979
timestamp 1649977179
transform 1 0 91172 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_981
timestamp 1649977179
transform 1 0 91356 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_993
timestamp 1649977179
transform 1 0 92460 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1005
timestamp 1649977179
transform 1 0 93564 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1017
timestamp 1649977179
transform 1 0 94668 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1029
timestamp 1649977179
transform 1 0 95772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1035
timestamp 1649977179
transform 1 0 96324 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1037
timestamp 1649977179
transform 1 0 96508 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1049
timestamp 1649977179
transform 1 0 97612 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1061
timestamp 1649977179
transform 1 0 98716 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1073
timestamp 1649977179
transform 1 0 99820 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1085
timestamp 1649977179
transform 1 0 100924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1091
timestamp 1649977179
transform 1 0 101476 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1093
timestamp 1649977179
transform 1 0 101660 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1105
timestamp 1649977179
transform 1 0 102764 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1117
timestamp 1649977179
transform 1 0 103868 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1129
timestamp 1649977179
transform 1 0 104972 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1141
timestamp 1649977179
transform 1 0 106076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1147
timestamp 1649977179
transform 1 0 106628 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1149
timestamp 1649977179
transform 1 0 106812 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1161
timestamp 1649977179
transform 1 0 107916 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1173
timestamp 1649977179
transform 1 0 109020 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1185
timestamp 1649977179
transform 1 0 110124 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1197
timestamp 1649977179
transform 1 0 111228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1203
timestamp 1649977179
transform 1 0 111780 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1205
timestamp 1649977179
transform 1 0 111964 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1217
timestamp 1649977179
transform 1 0 113068 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1229
timestamp 1649977179
transform 1 0 114172 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1241
timestamp 1649977179
transform 1 0 115276 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1253
timestamp 1649977179
transform 1 0 116380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1259
timestamp 1649977179
transform 1 0 116932 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1261
timestamp 1649977179
transform 1 0 117116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_1273
timestamp 1649977179
transform 1 0 118220 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_6
timestamp 1649977179
transform 1 0 1656 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_18
timestamp 1649977179
transform 1 0 2760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_30
timestamp 1649977179
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_42
timestamp 1649977179
transform 1 0 4968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1649977179
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1649977179
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1649977179
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1649977179
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1649977179
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1649977179
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1649977179
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1649977179
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1649977179
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1649977179
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1649977179
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1649977179
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_729
timestamp 1649977179
transform 1 0 68172 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_741
timestamp 1649977179
transform 1 0 69276 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_753
timestamp 1649977179
transform 1 0 70380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_765
timestamp 1649977179
transform 1 0 71484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 1649977179
transform 1 0 72588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 1649977179
transform 1 0 73140 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_785
timestamp 1649977179
transform 1 0 73324 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_797
timestamp 1649977179
transform 1 0 74428 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_809
timestamp 1649977179
transform 1 0 75532 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_821
timestamp 1649977179
transform 1 0 76636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_833
timestamp 1649977179
transform 1 0 77740 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_839
timestamp 1649977179
transform 1 0 78292 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_841
timestamp 1649977179
transform 1 0 78476 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_853
timestamp 1649977179
transform 1 0 79580 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_865
timestamp 1649977179
transform 1 0 80684 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_877
timestamp 1649977179
transform 1 0 81788 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_889
timestamp 1649977179
transform 1 0 82892 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_895
timestamp 1649977179
transform 1 0 83444 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_897
timestamp 1649977179
transform 1 0 83628 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_909
timestamp 1649977179
transform 1 0 84732 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_921
timestamp 1649977179
transform 1 0 85836 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_933
timestamp 1649977179
transform 1 0 86940 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_945
timestamp 1649977179
transform 1 0 88044 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_951
timestamp 1649977179
transform 1 0 88596 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_953
timestamp 1649977179
transform 1 0 88780 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_965
timestamp 1649977179
transform 1 0 89884 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_977
timestamp 1649977179
transform 1 0 90988 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_989
timestamp 1649977179
transform 1 0 92092 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1001
timestamp 1649977179
transform 1 0 93196 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1007
timestamp 1649977179
transform 1 0 93748 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1009
timestamp 1649977179
transform 1 0 93932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1021
timestamp 1649977179
transform 1 0 95036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1033
timestamp 1649977179
transform 1 0 96140 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1045
timestamp 1649977179
transform 1 0 97244 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1057
timestamp 1649977179
transform 1 0 98348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1063
timestamp 1649977179
transform 1 0 98900 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1065
timestamp 1649977179
transform 1 0 99084 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1077
timestamp 1649977179
transform 1 0 100188 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1089
timestamp 1649977179
transform 1 0 101292 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1101
timestamp 1649977179
transform 1 0 102396 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1113
timestamp 1649977179
transform 1 0 103500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1119
timestamp 1649977179
transform 1 0 104052 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1121
timestamp 1649977179
transform 1 0 104236 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1133
timestamp 1649977179
transform 1 0 105340 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1145
timestamp 1649977179
transform 1 0 106444 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1157
timestamp 1649977179
transform 1 0 107548 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1169
timestamp 1649977179
transform 1 0 108652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1175
timestamp 1649977179
transform 1 0 109204 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1177
timestamp 1649977179
transform 1 0 109388 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1189
timestamp 1649977179
transform 1 0 110492 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1201
timestamp 1649977179
transform 1 0 111596 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1213
timestamp 1649977179
transform 1 0 112700 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1225
timestamp 1649977179
transform 1 0 113804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1231
timestamp 1649977179
transform 1 0 114356 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1233
timestamp 1649977179
transform 1 0 114540 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1245
timestamp 1649977179
transform 1 0 115644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1257
timestamp 1649977179
transform 1 0 116748 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_1273
timestamp 1649977179
transform 1 0 118220 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_13
timestamp 1649977179
transform 1 0 2300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1649977179
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_319
timestamp 1649977179
transform 1 0 30452 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_330
timestamp 1649977179
transform 1 0 31464 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_342
timestamp 1649977179
transform 1 0 32568 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_354
timestamp 1649977179
transform 1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1649977179
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1649977179
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1649977179
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1649977179
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1649977179
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1649977179
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1649977179
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1649977179
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1649977179
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1649977179
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1649977179
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1649977179
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_725
timestamp 1649977179
transform 1 0 67804 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_737
timestamp 1649977179
transform 1 0 68908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 1649977179
transform 1 0 70012 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 1649977179
transform 1 0 70564 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_757
timestamp 1649977179
transform 1 0 70748 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_769
timestamp 1649977179
transform 1 0 71852 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_781
timestamp 1649977179
transform 1 0 72956 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_793
timestamp 1649977179
transform 1 0 74060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 1649977179
transform 1 0 75164 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 1649977179
transform 1 0 75716 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_813
timestamp 1649977179
transform 1 0 75900 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_825
timestamp 1649977179
transform 1 0 77004 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_837
timestamp 1649977179
transform 1 0 78108 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_849
timestamp 1649977179
transform 1 0 79212 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_861
timestamp 1649977179
transform 1 0 80316 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_867
timestamp 1649977179
transform 1 0 80868 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_869
timestamp 1649977179
transform 1 0 81052 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_881
timestamp 1649977179
transform 1 0 82156 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_893
timestamp 1649977179
transform 1 0 83260 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_905
timestamp 1649977179
transform 1 0 84364 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_917
timestamp 1649977179
transform 1 0 85468 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_923
timestamp 1649977179
transform 1 0 86020 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_925
timestamp 1649977179
transform 1 0 86204 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_937
timestamp 1649977179
transform 1 0 87308 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_949
timestamp 1649977179
transform 1 0 88412 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_961
timestamp 1649977179
transform 1 0 89516 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_973
timestamp 1649977179
transform 1 0 90620 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_979
timestamp 1649977179
transform 1 0 91172 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_981
timestamp 1649977179
transform 1 0 91356 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_993
timestamp 1649977179
transform 1 0 92460 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1005
timestamp 1649977179
transform 1 0 93564 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1017
timestamp 1649977179
transform 1 0 94668 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1029
timestamp 1649977179
transform 1 0 95772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1035
timestamp 1649977179
transform 1 0 96324 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1037
timestamp 1649977179
transform 1 0 96508 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1049
timestamp 1649977179
transform 1 0 97612 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1061
timestamp 1649977179
transform 1 0 98716 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1073
timestamp 1649977179
transform 1 0 99820 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1085
timestamp 1649977179
transform 1 0 100924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1091
timestamp 1649977179
transform 1 0 101476 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1093
timestamp 1649977179
transform 1 0 101660 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1105
timestamp 1649977179
transform 1 0 102764 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1117
timestamp 1649977179
transform 1 0 103868 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1129
timestamp 1649977179
transform 1 0 104972 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1141
timestamp 1649977179
transform 1 0 106076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1147
timestamp 1649977179
transform 1 0 106628 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1149
timestamp 1649977179
transform 1 0 106812 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1161
timestamp 1649977179
transform 1 0 107916 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1173
timestamp 1649977179
transform 1 0 109020 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1185
timestamp 1649977179
transform 1 0 110124 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1197
timestamp 1649977179
transform 1 0 111228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1203
timestamp 1649977179
transform 1 0 111780 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1205
timestamp 1649977179
transform 1 0 111964 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1217
timestamp 1649977179
transform 1 0 113068 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1229
timestamp 1649977179
transform 1 0 114172 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1241
timestamp 1649977179
transform 1 0 115276 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1253
timestamp 1649977179
transform 1 0 116380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1259
timestamp 1649977179
transform 1 0 116932 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1261
timestamp 1649977179
transform 1 0 117116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_1273
timestamp 1649977179
transform 1 0 118220 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_13
timestamp 1649977179
transform 1 0 2300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_25
timestamp 1649977179
transform 1 0 3404 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_37
timestamp 1649977179
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1649977179
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_330
timestamp 1649977179
transform 1 0 31464 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1649977179
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_346
timestamp 1649977179
transform 1 0 32936 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_350
timestamp 1649977179
transform 1 0 33304 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_362
timestamp 1649977179
transform 1 0 34408 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_374
timestamp 1649977179
transform 1 0 35512 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_386
timestamp 1649977179
transform 1 0 36616 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1649977179
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1649977179
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1649977179
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1649977179
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1649977179
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1649977179
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1649977179
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1649977179
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1649977179
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1649977179
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1649977179
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_729
timestamp 1649977179
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_741
timestamp 1649977179
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_753
timestamp 1649977179
transform 1 0 70380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_765
timestamp 1649977179
transform 1 0 71484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 1649977179
transform 1 0 72588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 1649977179
transform 1 0 73140 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_785
timestamp 1649977179
transform 1 0 73324 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_797
timestamp 1649977179
transform 1 0 74428 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_809
timestamp 1649977179
transform 1 0 75532 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_821
timestamp 1649977179
transform 1 0 76636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_833
timestamp 1649977179
transform 1 0 77740 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_839
timestamp 1649977179
transform 1 0 78292 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_841
timestamp 1649977179
transform 1 0 78476 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_853
timestamp 1649977179
transform 1 0 79580 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_865
timestamp 1649977179
transform 1 0 80684 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_877
timestamp 1649977179
transform 1 0 81788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_889
timestamp 1649977179
transform 1 0 82892 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_895
timestamp 1649977179
transform 1 0 83444 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_897
timestamp 1649977179
transform 1 0 83628 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_909
timestamp 1649977179
transform 1 0 84732 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_921
timestamp 1649977179
transform 1 0 85836 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_933
timestamp 1649977179
transform 1 0 86940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_945
timestamp 1649977179
transform 1 0 88044 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_951
timestamp 1649977179
transform 1 0 88596 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_953
timestamp 1649977179
transform 1 0 88780 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_965
timestamp 1649977179
transform 1 0 89884 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_977
timestamp 1649977179
transform 1 0 90988 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_989
timestamp 1649977179
transform 1 0 92092 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1001
timestamp 1649977179
transform 1 0 93196 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1007
timestamp 1649977179
transform 1 0 93748 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1009
timestamp 1649977179
transform 1 0 93932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1021
timestamp 1649977179
transform 1 0 95036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1033
timestamp 1649977179
transform 1 0 96140 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1045
timestamp 1649977179
transform 1 0 97244 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1057
timestamp 1649977179
transform 1 0 98348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1063
timestamp 1649977179
transform 1 0 98900 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1065
timestamp 1649977179
transform 1 0 99084 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1077
timestamp 1649977179
transform 1 0 100188 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1089
timestamp 1649977179
transform 1 0 101292 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1101
timestamp 1649977179
transform 1 0 102396 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1113
timestamp 1649977179
transform 1 0 103500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1119
timestamp 1649977179
transform 1 0 104052 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1121
timestamp 1649977179
transform 1 0 104236 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1133
timestamp 1649977179
transform 1 0 105340 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1145
timestamp 1649977179
transform 1 0 106444 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1157
timestamp 1649977179
transform 1 0 107548 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1169
timestamp 1649977179
transform 1 0 108652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1175
timestamp 1649977179
transform 1 0 109204 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1177
timestamp 1649977179
transform 1 0 109388 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1189
timestamp 1649977179
transform 1 0 110492 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1201
timestamp 1649977179
transform 1 0 111596 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1213
timestamp 1649977179
transform 1 0 112700 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1225
timestamp 1649977179
transform 1 0 113804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1231
timestamp 1649977179
transform 1 0 114356 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1233
timestamp 1649977179
transform 1 0 114540 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1245
timestamp 1649977179
transform 1 0 115644 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1257
timestamp 1649977179
transform 1 0 116748 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1265
timestamp 1649977179
transform 1 0 117484 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_1268
timestamp 1649977179
transform 1 0 117760 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_1273
timestamp 1649977179
transform 1 0 118220 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_341
timestamp 1649977179
transform 1 0 32476 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_346
timestamp 1649977179
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_358
timestamp 1649977179
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_481
timestamp 1649977179
transform 1 0 45356 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_493
timestamp 1649977179
transform 1 0 46460 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_505
timestamp 1649977179
transform 1 0 47564 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_517
timestamp 1649977179
transform 1 0 48668 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_529
timestamp 1649977179
transform 1 0 49772 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_620
timestamp 1649977179
transform 1 0 58144 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_632
timestamp 1649977179
transform 1 0 59248 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1649977179
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1649977179
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1649977179
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_681
timestamp 1649977179
transform 1 0 63756 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_687
timestamp 1649977179
transform 1 0 64308 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1649977179
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1649977179
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1649977179
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_725
timestamp 1649977179
transform 1 0 67804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_737
timestamp 1649977179
transform 1 0 68908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 1649977179
transform 1 0 70012 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 1649977179
transform 1 0 70564 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_757
timestamp 1649977179
transform 1 0 70748 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_769
timestamp 1649977179
transform 1 0 71852 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_781
timestamp 1649977179
transform 1 0 72956 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_793
timestamp 1649977179
transform 1 0 74060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 1649977179
transform 1 0 75164 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 1649977179
transform 1 0 75716 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_813
timestamp 1649977179
transform 1 0 75900 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_825
timestamp 1649977179
transform 1 0 77004 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_837
timestamp 1649977179
transform 1 0 78108 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_849
timestamp 1649977179
transform 1 0 79212 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_861
timestamp 1649977179
transform 1 0 80316 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_867
timestamp 1649977179
transform 1 0 80868 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_869
timestamp 1649977179
transform 1 0 81052 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_881
timestamp 1649977179
transform 1 0 82156 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_893
timestamp 1649977179
transform 1 0 83260 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_905
timestamp 1649977179
transform 1 0 84364 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_917
timestamp 1649977179
transform 1 0 85468 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_923
timestamp 1649977179
transform 1 0 86020 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_925
timestamp 1649977179
transform 1 0 86204 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_937
timestamp 1649977179
transform 1 0 87308 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_949
timestamp 1649977179
transform 1 0 88412 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_961
timestamp 1649977179
transform 1 0 89516 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_973
timestamp 1649977179
transform 1 0 90620 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_979
timestamp 1649977179
transform 1 0 91172 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_981
timestamp 1649977179
transform 1 0 91356 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_993
timestamp 1649977179
transform 1 0 92460 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1005
timestamp 1649977179
transform 1 0 93564 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1017
timestamp 1649977179
transform 1 0 94668 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1029
timestamp 1649977179
transform 1 0 95772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1035
timestamp 1649977179
transform 1 0 96324 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1037
timestamp 1649977179
transform 1 0 96508 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1049
timestamp 1649977179
transform 1 0 97612 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1061
timestamp 1649977179
transform 1 0 98716 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1073
timestamp 1649977179
transform 1 0 99820 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1085
timestamp 1649977179
transform 1 0 100924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1091
timestamp 1649977179
transform 1 0 101476 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1093
timestamp 1649977179
transform 1 0 101660 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1105
timestamp 1649977179
transform 1 0 102764 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1117
timestamp 1649977179
transform 1 0 103868 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1129
timestamp 1649977179
transform 1 0 104972 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1141
timestamp 1649977179
transform 1 0 106076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1147
timestamp 1649977179
transform 1 0 106628 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1149
timestamp 1649977179
transform 1 0 106812 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1161
timestamp 1649977179
transform 1 0 107916 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1173
timestamp 1649977179
transform 1 0 109020 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1185
timestamp 1649977179
transform 1 0 110124 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1197
timestamp 1649977179
transform 1 0 111228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1203
timestamp 1649977179
transform 1 0 111780 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1205
timestamp 1649977179
transform 1 0 111964 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1217
timestamp 1649977179
transform 1 0 113068 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1229
timestamp 1649977179
transform 1 0 114172 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1241
timestamp 1649977179
transform 1 0 115276 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1253
timestamp 1649977179
transform 1 0 116380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1259
timestamp 1649977179
transform 1 0 116932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_1261
timestamp 1649977179
transform 1 0 117116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1269
timestamp 1649977179
transform 1 0 117852 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_1273
timestamp 1649977179
transform 1 0 118220 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_6
timestamp 1649977179
transform 1 0 1656 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_18
timestamp 1649977179
transform 1 0 2760 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_30
timestamp 1649977179
transform 1 0 3864 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_42
timestamp 1649977179
transform 1 0 4968 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1649977179
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_369
timestamp 1649977179
transform 1 0 35052 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_374
timestamp 1649977179
transform 1 0 35512 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_386
timestamp 1649977179
transform 1 0 36616 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_622
timestamp 1649977179
transform 1 0 58328 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_626
timestamp 1649977179
transform 1 0 58696 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_634
timestamp 1649977179
transform 1 0 59432 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_637
timestamp 1649977179
transform 1 0 59708 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_648
timestamp 1649977179
transform 1 0 60720 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_656
timestamp 1649977179
transform 1 0 61456 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_661
timestamp 1649977179
transform 1 0 61916 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_669
timestamp 1649977179
transform 1 0 62652 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1649977179
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1649977179
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1649977179
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1649977179
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1649977179
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1649977179
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_729
timestamp 1649977179
transform 1 0 68172 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_741
timestamp 1649977179
transform 1 0 69276 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_753
timestamp 1649977179
transform 1 0 70380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_765
timestamp 1649977179
transform 1 0 71484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 1649977179
transform 1 0 72588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 1649977179
transform 1 0 73140 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_785
timestamp 1649977179
transform 1 0 73324 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_797
timestamp 1649977179
transform 1 0 74428 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_809
timestamp 1649977179
transform 1 0 75532 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_818
timestamp 1649977179
transform 1 0 76360 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_830
timestamp 1649977179
transform 1 0 77464 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_838
timestamp 1649977179
transform 1 0 78200 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_841
timestamp 1649977179
transform 1 0 78476 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_853
timestamp 1649977179
transform 1 0 79580 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_865
timestamp 1649977179
transform 1 0 80684 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_877
timestamp 1649977179
transform 1 0 81788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_889
timestamp 1649977179
transform 1 0 82892 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_895
timestamp 1649977179
transform 1 0 83444 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_897
timestamp 1649977179
transform 1 0 83628 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_909
timestamp 1649977179
transform 1 0 84732 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_921
timestamp 1649977179
transform 1 0 85836 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_933
timestamp 1649977179
transform 1 0 86940 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_945
timestamp 1649977179
transform 1 0 88044 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_951
timestamp 1649977179
transform 1 0 88596 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_953
timestamp 1649977179
transform 1 0 88780 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_965
timestamp 1649977179
transform 1 0 89884 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_977
timestamp 1649977179
transform 1 0 90988 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_989
timestamp 1649977179
transform 1 0 92092 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1001
timestamp 1649977179
transform 1 0 93196 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1007
timestamp 1649977179
transform 1 0 93748 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1009
timestamp 1649977179
transform 1 0 93932 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1021
timestamp 1649977179
transform 1 0 95036 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1033
timestamp 1649977179
transform 1 0 96140 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1045
timestamp 1649977179
transform 1 0 97244 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1057
timestamp 1649977179
transform 1 0 98348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1063
timestamp 1649977179
transform 1 0 98900 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1065
timestamp 1649977179
transform 1 0 99084 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1077
timestamp 1649977179
transform 1 0 100188 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1089
timestamp 1649977179
transform 1 0 101292 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1101
timestamp 1649977179
transform 1 0 102396 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1113
timestamp 1649977179
transform 1 0 103500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1119
timestamp 1649977179
transform 1 0 104052 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1121
timestamp 1649977179
transform 1 0 104236 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1133
timestamp 1649977179
transform 1 0 105340 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1145
timestamp 1649977179
transform 1 0 106444 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1157
timestamp 1649977179
transform 1 0 107548 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1169
timestamp 1649977179
transform 1 0 108652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1175
timestamp 1649977179
transform 1 0 109204 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1177
timestamp 1649977179
transform 1 0 109388 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1189
timestamp 1649977179
transform 1 0 110492 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1201
timestamp 1649977179
transform 1 0 111596 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1213
timestamp 1649977179
transform 1 0 112700 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1225
timestamp 1649977179
transform 1 0 113804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1231
timestamp 1649977179
transform 1 0 114356 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1233
timestamp 1649977179
transform 1 0 114540 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1245
timestamp 1649977179
transform 1 0 115644 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_1257
timestamp 1649977179
transform 1 0 116748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1261
timestamp 1649977179
transform 1 0 117116 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_1265
timestamp 1649977179
transform 1 0 117484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_1273
timestamp 1649977179
transform 1 0 118220 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_13
timestamp 1649977179
transform 1 0 2300 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1649977179
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_314
timestamp 1649977179
transform 1 0 29992 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_326
timestamp 1649977179
transform 1 0 31096 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_338
timestamp 1649977179
transform 1 0 32200 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_350
timestamp 1649977179
transform 1 0 33304 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1649977179
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_369
timestamp 1649977179
transform 1 0 35052 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_379
timestamp 1649977179
transform 1 0 35972 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_391
timestamp 1649977179
transform 1 0 37076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_403
timestamp 1649977179
transform 1 0 38180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_415
timestamp 1649977179
transform 1 0 39284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_496
timestamp 1649977179
transform 1 0 46736 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_508
timestamp 1649977179
transform 1 0 47840 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_524
timestamp 1649977179
transform 1 0 49312 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_536
timestamp 1649977179
transform 1 0 50416 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_548
timestamp 1649977179
transform 1 0 51520 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_560
timestamp 1649977179
transform 1 0 52624 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_568
timestamp 1649977179
transform 1 0 53360 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_573
timestamp 1649977179
transform 1 0 53820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_584
timestamp 1649977179
transform 1 0 54832 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_592
timestamp 1649977179
transform 1 0 55568 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_600
timestamp 1649977179
transform 1 0 56304 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_604
timestamp 1649977179
transform 1 0 56672 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_616
timestamp 1649977179
transform 1 0 57776 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_624
timestamp 1649977179
transform 1 0 58512 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_629
timestamp 1649977179
transform 1 0 58972 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_641
timestamp 1649977179
transform 1 0 60076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_645
timestamp 1649977179
transform 1 0 60444 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_653
timestamp 1649977179
transform 1 0 61180 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_663
timestamp 1649977179
transform 1 0 62100 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_670
timestamp 1649977179
transform 1 0 62744 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_682
timestamp 1649977179
transform 1 0 63848 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_694
timestamp 1649977179
transform 1 0 64952 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1649977179
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1649977179
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_725
timestamp 1649977179
transform 1 0 67804 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_737
timestamp 1649977179
transform 1 0 68908 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_742
timestamp 1649977179
transform 1 0 69368 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_748
timestamp 1649977179
transform 1 0 69920 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_752
timestamp 1649977179
transform 1 0 70288 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_757
timestamp 1649977179
transform 1 0 70748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_765
timestamp 1649977179
transform 1 0 71484 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_772
timestamp 1649977179
transform 1 0 72128 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_784
timestamp 1649977179
transform 1 0 73232 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_796
timestamp 1649977179
transform 1 0 74336 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_800
timestamp 1649977179
transform 1 0 74704 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_804
timestamp 1649977179
transform 1 0 75072 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_813
timestamp 1649977179
transform 1 0 75900 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_823
timestamp 1649977179
transform 1 0 76820 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_832
timestamp 1649977179
transform 1 0 77648 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_844
timestamp 1649977179
transform 1 0 78752 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_857
timestamp 1649977179
transform 1 0 79948 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_865
timestamp 1649977179
transform 1 0 80684 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_869
timestamp 1649977179
transform 1 0 81052 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_881
timestamp 1649977179
transform 1 0 82156 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_893
timestamp 1649977179
transform 1 0 83260 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_905
timestamp 1649977179
transform 1 0 84364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_917
timestamp 1649977179
transform 1 0 85468 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_923
timestamp 1649977179
transform 1 0 86020 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_925
timestamp 1649977179
transform 1 0 86204 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_937
timestamp 1649977179
transform 1 0 87308 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_949
timestamp 1649977179
transform 1 0 88412 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_961
timestamp 1649977179
transform 1 0 89516 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_972
timestamp 1649977179
transform 1 0 90528 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_981
timestamp 1649977179
transform 1 0 91356 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_989
timestamp 1649977179
transform 1 0 92092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_1001
timestamp 1649977179
transform 1 0 93196 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1007
timestamp 1649977179
transform 1 0 93748 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1019
timestamp 1649977179
transform 1 0 94852 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_1031
timestamp 1649977179
transform 1 0 95956 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1035
timestamp 1649977179
transform 1 0 96324 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1037
timestamp 1649977179
transform 1 0 96508 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1049
timestamp 1649977179
transform 1 0 97612 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1061
timestamp 1649977179
transform 1 0 98716 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1073
timestamp 1649977179
transform 1 0 99820 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1085
timestamp 1649977179
transform 1 0 100924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1091
timestamp 1649977179
transform 1 0 101476 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1093
timestamp 1649977179
transform 1 0 101660 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1105
timestamp 1649977179
transform 1 0 102764 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1117
timestamp 1649977179
transform 1 0 103868 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1129
timestamp 1649977179
transform 1 0 104972 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1141
timestamp 1649977179
transform 1 0 106076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1147
timestamp 1649977179
transform 1 0 106628 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1149
timestamp 1649977179
transform 1 0 106812 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1161
timestamp 1649977179
transform 1 0 107916 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1173
timestamp 1649977179
transform 1 0 109020 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1185
timestamp 1649977179
transform 1 0 110124 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1197
timestamp 1649977179
transform 1 0 111228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1203
timestamp 1649977179
transform 1 0 111780 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1205
timestamp 1649977179
transform 1 0 111964 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1217
timestamp 1649977179
transform 1 0 113068 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1229
timestamp 1649977179
transform 1 0 114172 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1241
timestamp 1649977179
transform 1 0 115276 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1253
timestamp 1649977179
transform 1 0 116380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1259
timestamp 1649977179
transform 1 0 116932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_1265
timestamp 1649977179
transform 1 0 117484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_1273
timestamp 1649977179
transform 1 0 118220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_13
timestamp 1649977179
transform 1 0 2300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_20
timestamp 1649977179
transform 1 0 2944 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_35
timestamp 1649977179
transform 1 0 4324 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_41
timestamp 1649977179
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1649977179
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_76
timestamp 1649977179
transform 1 0 8096 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_88
timestamp 1649977179
transform 1 0 9200 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_100
timestamp 1649977179
transform 1 0 10304 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_106
timestamp 1649977179
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_118
timestamp 1649977179
transform 1 0 11960 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_130
timestamp 1649977179
transform 1 0 13064 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_142
timestamp 1649977179
transform 1 0 14168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_153
timestamp 1649977179
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_201
timestamp 1649977179
transform 1 0 19596 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_207
timestamp 1649977179
transform 1 0 20148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_214
timestamp 1649977179
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1649977179
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_286
timestamp 1649977179
transform 1 0 27416 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_298
timestamp 1649977179
transform 1 0 28520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_306
timestamp 1649977179
transform 1 0 29256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_310
timestamp 1649977179
transform 1 0 29624 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_323
timestamp 1649977179
transform 1 0 30820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_345
timestamp 1649977179
transform 1 0 32844 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_355
timestamp 1649977179
transform 1 0 33764 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_359
timestamp 1649977179
transform 1 0 34132 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_367
timestamp 1649977179
transform 1 0 34868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_380
timestamp 1649977179
transform 1 0 36064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 1649977179
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_401
timestamp 1649977179
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_413
timestamp 1649977179
transform 1 0 39100 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_424
timestamp 1649977179
transform 1 0 40112 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_431
timestamp 1649977179
transform 1 0 40756 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_440
timestamp 1649977179
transform 1 0 41584 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_489
timestamp 1649977179
transform 1 0 46092 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_493
timestamp 1649977179
transform 1 0 46460 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_500
timestamp 1649977179
transform 1 0 47104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_509
timestamp 1649977179
transform 1 0 47932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_520
timestamp 1649977179
transform 1 0 48944 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_527
timestamp 1649977179
transform 1 0 49588 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_534
timestamp 1649977179
transform 1 0 50232 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_542
timestamp 1649977179
transform 1 0 50968 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_550
timestamp 1649977179
transform 1 0 51704 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_558
timestamp 1649977179
transform 1 0 52440 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_566
timestamp 1649977179
transform 1 0 53176 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_581
timestamp 1649977179
transform 1 0 54556 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_601
timestamp 1649977179
transform 1 0 56396 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_605
timestamp 1649977179
transform 1 0 56764 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_612
timestamp 1649977179
transform 1 0 57408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_623
timestamp 1649977179
transform 1 0 58420 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_636
timestamp 1649977179
transform 1 0 59616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_650
timestamp 1649977179
transform 1 0 60904 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_656
timestamp 1649977179
transform 1 0 61456 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_666
timestamp 1649977179
transform 1 0 62376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_670
timestamp 1649977179
transform 1 0 62744 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_673
timestamp 1649977179
transform 1 0 63020 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_685
timestamp 1649977179
transform 1 0 64124 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_698
timestamp 1649977179
transform 1 0 65320 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_705
timestamp 1649977179
transform 1 0 65964 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_712
timestamp 1649977179
transform 1 0 66608 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_724
timestamp 1649977179
transform 1 0 67712 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1649977179
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_739
timestamp 1649977179
transform 1 0 69092 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_747
timestamp 1649977179
transform 1 0 69828 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_753
timestamp 1649977179
transform 1 0 70380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_760
timestamp 1649977179
transform 1 0 71024 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_768
timestamp 1649977179
transform 1 0 71760 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_778
timestamp 1649977179
transform 1 0 72680 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_805
timestamp 1649977179
transform 1 0 75164 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_809
timestamp 1649977179
transform 1 0 75532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_819
timestamp 1649977179
transform 1 0 76452 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_823
timestamp 1649977179
transform 1 0 76820 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_834
timestamp 1649977179
transform 1 0 77832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_838
timestamp 1649977179
transform 1 0 78200 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_844
timestamp 1649977179
transform 1 0 78752 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_851
timestamp 1649977179
transform 1 0 79396 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_858
timestamp 1649977179
transform 1 0 80040 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_870
timestamp 1649977179
transform 1 0 81144 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_882
timestamp 1649977179
transform 1 0 82248 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_894
timestamp 1649977179
transform 1 0 83352 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_897
timestamp 1649977179
transform 1 0 83628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_905
timestamp 1649977179
transform 1 0 84364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_912
timestamp 1649977179
transform 1 0 85008 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_919
timestamp 1649977179
transform 1 0 85652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_926
timestamp 1649977179
transform 1 0 86296 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_933
timestamp 1649977179
transform 1 0 86940 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_945
timestamp 1649977179
transform 1 0 88044 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_951
timestamp 1649977179
transform 1 0 88596 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_953
timestamp 1649977179
transform 1 0 88780 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_959
timestamp 1649977179
transform 1 0 89332 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_963
timestamp 1649977179
transform 1 0 89700 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_974
timestamp 1649977179
transform 1 0 90712 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_978
timestamp 1649977179
transform 1 0 91080 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_986
timestamp 1649977179
transform 1 0 91816 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_993
timestamp 1649977179
transform 1 0 92460 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1000
timestamp 1649977179
transform 1 0 93104 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1009
timestamp 1649977179
transform 1 0 93932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1017
timestamp 1649977179
transform 1 0 94668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1024
timestamp 1649977179
transform 1 0 95312 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1031
timestamp 1649977179
transform 1 0 95956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1043
timestamp 1649977179
transform 1 0 97060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1055
timestamp 1649977179
transform 1 0 98164 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1063
timestamp 1649977179
transform 1 0 98900 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1065
timestamp 1649977179
transform 1 0 99084 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1077
timestamp 1649977179
transform 1 0 100188 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1084
timestamp 1649977179
transform 1 0 100832 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1096
timestamp 1649977179
transform 1 0 101936 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1108
timestamp 1649977179
transform 1 0 103040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1112
timestamp 1649977179
transform 1 0 103408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1116
timestamp 1649977179
transform 1 0 103776 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1121
timestamp 1649977179
transform 1 0 104236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1129
timestamp 1649977179
transform 1 0 104972 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1136
timestamp 1649977179
transform 1 0 105616 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1148
timestamp 1649977179
transform 1 0 106720 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1160
timestamp 1649977179
transform 1 0 107824 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1172
timestamp 1649977179
transform 1 0 108928 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1177
timestamp 1649977179
transform 1 0 109388 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1189
timestamp 1649977179
transform 1 0 110492 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_1197
timestamp 1649977179
transform 1 0 111228 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1203
timestamp 1649977179
transform 1 0 111780 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1215
timestamp 1649977179
transform 1 0 112884 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1227
timestamp 1649977179
transform 1 0 113988 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1231
timestamp 1649977179
transform 1 0 114356 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1233
timestamp 1649977179
transform 1 0 114540 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1245
timestamp 1649977179
transform 1 0 115644 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1251
timestamp 1649977179
transform 1 0 116196 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_1255
timestamp 1649977179
transform 1 0 116564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_1259
timestamp 1649977179
transform 1 0 116932 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_1265
timestamp 1649977179
transform 1 0 117484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1273
timestamp 1649977179
transform 1 0 118220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_6
timestamp 1649977179
transform 1 0 1656 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1649977179
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_37
timestamp 1649977179
transform 1 0 4508 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_52
timestamp 1649977179
transform 1 0 5888 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_67
timestamp 1649977179
transform 1 0 7268 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_71
timestamp 1649977179
transform 1 0 7636 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_95
timestamp 1649977179
transform 1 0 9844 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_103
timestamp 1649977179
transform 1 0 10580 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_107
timestamp 1649977179
transform 1 0 10948 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_110
timestamp 1649977179
transform 1 0 11224 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_117
timestamp 1649977179
transform 1 0 11868 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_126
timestamp 1649977179
transform 1 0 12696 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1649977179
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_144
timestamp 1649977179
transform 1 0 14352 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_152
timestamp 1649977179
transform 1 0 15088 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_164
timestamp 1649977179
transform 1 0 16192 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_169
timestamp 1649977179
transform 1 0 16652 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_173
timestamp 1649977179
transform 1 0 17020 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_178
timestamp 1649977179
transform 1 0 17480 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1649977179
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_200
timestamp 1649977179
transform 1 0 19504 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_210
timestamp 1649977179
transform 1 0 20424 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_217
timestamp 1649977179
transform 1 0 21068 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_223
timestamp 1649977179
transform 1 0 21620 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_225
timestamp 1649977179
transform 1 0 21804 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_230
timestamp 1649977179
transform 1 0 22264 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_237
timestamp 1649977179
transform 1 0 22908 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1649977179
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_256
timestamp 1649977179
transform 1 0 24656 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_260
timestamp 1649977179
transform 1 0 25024 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_266
timestamp 1649977179
transform 1 0 25576 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_270
timestamp 1649977179
transform 1 0 25944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_278
timestamp 1649977179
transform 1 0 26680 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_285
timestamp 1649977179
transform 1 0 27324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_294
timestamp 1649977179
transform 1 0 28152 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_298
timestamp 1649977179
transform 1 0 28520 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1649977179
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_324
timestamp 1649977179
transform 1 0 30912 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_332
timestamp 1649977179
transform 1 0 31648 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_337
timestamp 1649977179
transform 1 0 32108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_349
timestamp 1649977179
transform 1 0 33212 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1649977179
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_375
timestamp 1649977179
transform 1 0 35604 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_379
timestamp 1649977179
transform 1 0 35972 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_385
timestamp 1649977179
transform 1 0 36524 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_393
timestamp 1649977179
transform 1 0 37260 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_405
timestamp 1649977179
transform 1 0 38364 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_409
timestamp 1649977179
transform 1 0 38732 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_416
timestamp 1649977179
transform 1 0 39376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_430
timestamp 1649977179
transform 1 0 40664 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_434
timestamp 1649977179
transform 1 0 41032 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_444
timestamp 1649977179
transform 1 0 41952 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_453
timestamp 1649977179
transform 1 0 42780 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_460
timestamp 1649977179
transform 1 0 43424 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_464
timestamp 1649977179
transform 1 0 43792 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_468
timestamp 1649977179
transform 1 0 44160 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_480
timestamp 1649977179
transform 1 0 45264 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_486
timestamp 1649977179
transform 1 0 45816 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_491
timestamp 1649977179
transform 1 0 46276 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_500
timestamp 1649977179
transform 1 0 47104 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_505
timestamp 1649977179
transform 1 0 47564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_509
timestamp 1649977179
transform 1 0 47932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_514
timestamp 1649977179
transform 1 0 48392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_527
timestamp 1649977179
transform 1 0 49588 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_538
timestamp 1649977179
transform 1 0 50600 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_556
timestamp 1649977179
transform 1 0 52256 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_561
timestamp 1649977179
transform 1 0 52716 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_567
timestamp 1649977179
transform 1 0 53268 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_571
timestamp 1649977179
transform 1 0 53636 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_582
timestamp 1649977179
transform 1 0 54648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_586
timestamp 1649977179
transform 1 0 55016 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_593
timestamp 1649977179
transform 1 0 55660 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_599
timestamp 1649977179
transform 1 0 56212 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_602
timestamp 1649977179
transform 1 0 56488 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_612
timestamp 1649977179
transform 1 0 57408 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_617
timestamp 1649977179
transform 1 0 57868 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_621
timestamp 1649977179
transform 1 0 58236 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_632
timestamp 1649977179
transform 1 0 59248 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_639
timestamp 1649977179
transform 1 0 59892 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1649977179
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_645
timestamp 1649977179
transform 1 0 60444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_656
timestamp 1649977179
transform 1 0 61456 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_663
timestamp 1649977179
transform 1 0 62100 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_671
timestamp 1649977179
transform 1 0 62836 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_673
timestamp 1649977179
transform 1 0 63020 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_685
timestamp 1649977179
transform 1 0 64124 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_692
timestamp 1649977179
transform 1 0 64768 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_704
timestamp 1649977179
transform 1 0 65872 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_711
timestamp 1649977179
transform 1 0 66516 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_718
timestamp 1649977179
transform 1 0 67160 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_726
timestamp 1649977179
transform 1 0 67896 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_738
timestamp 1649977179
transform 1 0 69000 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_745
timestamp 1649977179
transform 1 0 69644 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_752
timestamp 1649977179
transform 1 0 70288 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_766
timestamp 1649977179
transform 1 0 71576 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_780
timestamp 1649977179
transform 1 0 72864 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_785
timestamp 1649977179
transform 1 0 73324 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_793
timestamp 1649977179
transform 1 0 74060 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_797
timestamp 1649977179
transform 1 0 74428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_808
timestamp 1649977179
transform 1 0 75440 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_816
timestamp 1649977179
transform 1 0 76176 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_832
timestamp 1649977179
transform 1 0 77648 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_841
timestamp 1649977179
transform 1 0 78476 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_852
timestamp 1649977179
transform 1 0 79488 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_859
timestamp 1649977179
transform 1 0 80132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_867
timestamp 1649977179
transform 1 0 80868 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_873
timestamp 1649977179
transform 1 0 81420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_880
timestamp 1649977179
transform 1 0 82064 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_884
timestamp 1649977179
transform 1 0 82432 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_888
timestamp 1649977179
transform 1 0 82800 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_900
timestamp 1649977179
transform 1 0 83904 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_915
timestamp 1649977179
transform 1 0 85284 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_923
timestamp 1649977179
transform 1 0 86020 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_928
timestamp 1649977179
transform 1 0 86480 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_937
timestamp 1649977179
transform 1 0 87308 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_944
timestamp 1649977179
transform 1 0 87952 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_956
timestamp 1649977179
transform 1 0 89056 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_961
timestamp 1649977179
transform 1 0 89516 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_965
timestamp 1649977179
transform 1 0 89884 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_976
timestamp 1649977179
transform 1 0 90896 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_981
timestamp 1649977179
transform 1 0 91356 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_991
timestamp 1649977179
transform 1 0 92276 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_999
timestamp 1649977179
transform 1 0 93012 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1007
timestamp 1649977179
transform 1 0 93748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1009
timestamp 1649977179
transform 1 0 93932 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1022
timestamp 1649977179
transform 1 0 95128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1029
timestamp 1649977179
transform 1 0 95772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1035
timestamp 1649977179
transform 1 0 96324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1040
timestamp 1649977179
transform 1 0 96784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1047
timestamp 1649977179
transform 1 0 97428 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1056
timestamp 1649977179
transform 1 0 98256 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1075
timestamp 1649977179
transform 1 0 100004 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1082
timestamp 1649977179
transform 1 0 100648 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_1090
timestamp 1649977179
transform 1 0 101384 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1096
timestamp 1649977179
transform 1 0 101936 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1105
timestamp 1649977179
transform 1 0 102764 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1112
timestamp 1649977179
transform 1 0 103408 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1121
timestamp 1649977179
transform 1 0 104236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1129
timestamp 1649977179
transform 1 0 104972 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1137
timestamp 1649977179
transform 1 0 105708 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1144
timestamp 1649977179
transform 1 0 106352 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1149
timestamp 1649977179
transform 1 0 106812 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_1157
timestamp 1649977179
transform 1 0 107548 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_1161
timestamp 1649977179
transform 1 0 107916 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1168
timestamp 1649977179
transform 1 0 108560 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1180
timestamp 1649977179
transform 1 0 109664 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1187
timestamp 1649977179
transform 1 0 110308 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1196
timestamp 1649977179
transform 1 0 111136 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1205
timestamp 1649977179
transform 1 0 111964 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1213
timestamp 1649977179
transform 1 0 112700 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1224
timestamp 1649977179
transform 1 0 113712 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1236
timestamp 1649977179
transform 1 0 114816 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1245
timestamp 1649977179
transform 1 0 115644 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1253
timestamp 1649977179
transform 1 0 116380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1259
timestamp 1649977179
transform 1 0 116932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_1261
timestamp 1649977179
transform 1 0 117116 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1273
timestamp 1649977179
transform 1 0 118220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 118864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 118864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 118864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 118864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 118864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 118864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 118864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 118864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 118864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 118864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 118864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 118864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 118864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 118864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 118864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 118864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 118864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 118864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 118864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 118864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 118864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 118864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 118864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 118864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 118864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 118864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 118864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 118864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 118864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 118864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 118864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 118864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 118864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 118864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 118864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 118864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 118864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 118864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 118864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 118864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 118864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 118864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 118864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 118864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 118864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 118864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 118864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 80960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 86112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 91264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 96416 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 101568 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 106720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 111872 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 117024 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 83536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 88688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 93840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 98992 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 104144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 109296 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 114448 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 80960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 86112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 91264 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 96416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 101568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 106720 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 111872 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 117024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 83536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 88688 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 93840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 98992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 104144 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 109296 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 114448 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 80960 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 86112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 91264 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 96416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 101568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 106720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 111872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 117024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 83536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 88688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 93840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 98992 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 104144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 109296 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 114448 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 80960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 86112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 91264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 96416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 101568 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 106720 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 111872 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 117024 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 83536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 88688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 93840 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 98992 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 104144 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 109296 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 114448 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 80960 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 86112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 91264 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 96416 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 101568 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 106720 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 111872 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 117024 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 83536 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 88688 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 93840 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 98992 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 104144 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 109296 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 114448 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 80960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 86112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 91264 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 96416 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 101568 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 106720 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 111872 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 117024 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 83536 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 88688 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 93840 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 98992 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 104144 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 109296 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 114448 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 80960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 86112 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 91264 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 96416 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 101568 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 106720 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 111872 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 117024 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 83536 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 88688 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 93840 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 98992 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 104144 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 109296 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 114448 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 70656 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 75808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 80960 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 86112 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 91264 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 96416 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 101568 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 106720 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 111872 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 117024 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 73232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 78384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 83536 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 88688 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 93840 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 98992 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 104144 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 109296 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 114448 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 70656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 75808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 80960 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 86112 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 91264 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 96416 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 101568 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 106720 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 111872 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 117024 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 73232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 78384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 83536 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 88688 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 93840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 98992 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 104144 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 109296 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 114448 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 70656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 75808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 80960 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 86112 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 91264 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 96416 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 101568 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 106720 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 111872 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 117024 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 73232 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 78384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 83536 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 88688 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 93840 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 98992 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 104144 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 109296 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 114448 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 70656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 75808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 80960 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 86112 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 91264 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 96416 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 101568 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 106720 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 111872 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 117024 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 73232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 78384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 83536 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 88688 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 93840 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 98992 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 104144 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 109296 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 114448 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 70656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 75808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 80960 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 86112 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 91264 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 96416 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 101568 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 106720 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 111872 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 117024 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 73232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 78384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 83536 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 88688 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 93840 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 98992 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 104144 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 109296 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 114448 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 70656 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 75808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 80960 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 86112 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 91264 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 96416 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 101568 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 106720 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 111872 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 117024 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 73232 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 78384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 83536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 88688 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 93840 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 98992 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 104144 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 109296 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 114448 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 70656 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 75808 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 80960 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 86112 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 91264 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 96416 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 101568 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 106720 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 111872 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 117024 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 73232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 78384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 83536 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 88688 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 93840 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 98992 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 104144 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 109296 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 114448 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 70656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 75808 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 80960 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 86112 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 91264 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 96416 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 101568 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 106720 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 111872 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 117024 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 73232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 78384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 83536 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 88688 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 93840 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 98992 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 104144 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 109296 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 114448 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 70656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 75808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 80960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 86112 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 91264 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 96416 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 101568 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 106720 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 111872 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 117024 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 73232 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 78384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 83536 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 88688 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 93840 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 98992 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 104144 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 109296 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 114448 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 32016 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 37168 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 42320 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 47472 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 52624 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 57776 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 62928 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 68080 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 70656 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 73232 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 75808 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 78384 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 80960 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 83536 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 86112 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 88688 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 91264 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 93840 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 96416 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 98992 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 101568 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 104144 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 106720 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 109296 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 111872 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 114448 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 117024 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _106_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 69184 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _107_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 69276 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _108_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 70748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _109_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 68080 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _110_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 69460 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _111_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 70748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _112_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 71484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _113_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 70748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _114_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 67988 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _115_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 67068 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _116_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 66792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1649977179
transform 1 0 70012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _118_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 69920 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _119_
timestamp 1649977179
transform 1 0 68172 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _120_
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _121_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 66884 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1649977179
transform 1 0 64676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _123_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 65780 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _124_
timestamp 1649977179
transform 1 0 84456 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _125_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 83628 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _126_
timestamp 1649977179
transform 1 0 56580 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1649977179
transform 1 0 55752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _128_
timestamp 1649977179
transform 1 0 84456 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1649977179
transform 1 0 86020 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _131_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43700 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _132_
timestamp 1649977179
transform 1 0 76360 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1649977179
transform 1 0 76820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 1649977179
transform 1 0 76544 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1649977179
transform 1 0 74428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _136_
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1649977179
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _138_
timestamp 1649977179
transform 1 0 29716 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _139_
timestamp 1649977179
transform 1 0 29440 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _140_
timestamp 1649977179
transform 1 0 76452 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1649977179
transform 1 0 76912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _142_
timestamp 1649977179
transform 1 0 54464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _143_
timestamp 1649977179
transform 1 0 55292 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _144_
timestamp 1649977179
transform 1 0 53636 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _145_
timestamp 1649977179
transform 1 0 77004 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1649977179
transform 1 0 78476 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _147_
timestamp 1649977179
transform 1 0 72312 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _148_
timestamp 1649977179
transform 1 0 71852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _149_
timestamp 1649977179
transform 1 0 75624 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _150_
timestamp 1649977179
transform 1 0 76452 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _151_
timestamp 1649977179
transform 1 0 68172 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _152_
timestamp 1649977179
transform 1 0 68540 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _153_
timestamp 1649977179
transform 1 0 55660 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _154_
timestamp 1649977179
transform 1 0 78660 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1649977179
transform 1 0 79212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _156_
timestamp 1649977179
transform 1 0 68172 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1649977179
transform 1 0 68448 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _158_
timestamp 1649977179
transform 1 0 78660 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1649977179
transform 1 0 79948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _160_
timestamp 1649977179
transform 1 0 74612 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _161_
timestamp 1649977179
transform 1 0 74244 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _162_
timestamp 1649977179
transform 1 0 53820 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1649977179
transform 1 0 53268 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _164_
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _165_
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1649977179
transform 1 0 49220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _167_
timestamp 1649977179
transform 1 0 48760 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1649977179
transform 1 0 49312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _169_
timestamp 1649977179
transform 1 0 35144 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _170_
timestamp 1649977179
transform 1 0 48024 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _171_
timestamp 1649977179
transform 1 0 35236 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1649977179
transform 1 0 33856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _173_
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp 1649977179
transform 1 0 40480 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _175_
timestamp 1649977179
transform 1 0 54556 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _176_
timestamp 1649977179
transform 1 0 50508 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _177_
timestamp 1649977179
transform 1 0 58788 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _178_
timestamp 1649977179
transform 1 0 59432 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _179_
timestamp 1649977179
transform 1 0 70748 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _180_
timestamp 1649977179
transform 1 0 71116 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _181_
timestamp 1649977179
transform 1 0 42596 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _182_
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _183_
timestamp 1649977179
transform 1 0 52716 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1649977179
transform 1 0 51796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1649977179
transform 1 0 69276 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1649977179
transform 1 0 70288 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _187_
timestamp 1649977179
transform 1 0 55844 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _188_
timestamp 1649977179
transform 1 0 70748 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp 1649977179
transform 1 0 70748 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _190_
timestamp 1649977179
transform 1 0 29992 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _191_
timestamp 1649977179
transform 1 0 39192 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _192_
timestamp 1649977179
transform 1 0 85836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1649977179
transform 1 0 86572 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _194_
timestamp 1649977179
transform 1 0 30084 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1649977179
transform 1 0 29348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp 1649977179
transform 1 0 61548 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1649977179
transform 1 0 61640 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _198_
timestamp 1649977179
transform 1 0 53636 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _199_
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _200_
timestamp 1649977179
transform 1 0 41492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp 1649977179
transform 1 0 65596 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1649977179
transform 1 0 65596 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp 1649977179
transform 1 0 51428 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1649977179
transform 1 0 50784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1649977179
transform 1 0 66148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 1649977179
transform 1 0 40020 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _208_
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _209_
timestamp 1649977179
transform 1 0 49496 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 1649977179
transform 1 0 33304 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _211_
timestamp 1649977179
transform 1 0 33028 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1649977179
transform 1 0 38088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 1649977179
transform 1 0 35972 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _215_
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _217_
timestamp 1649977179
transform 1 0 36524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1649977179
transform 1 0 30636 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1649977179
transform 1 0 45080 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _220_
timestamp 1649977179
transform 1 0 50416 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 1649977179
transform 1 0 22080 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _223_
timestamp 1649977179
transform 1 0 38824 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _224_
timestamp 1649977179
transform 1 0 42504 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 1649977179
transform 1 0 64492 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1649977179
transform 1 0 65688 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _227_
timestamp 1649977179
transform 1 0 63296 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _228_
timestamp 1649977179
transform 1 0 63940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _229_
timestamp 1649977179
transform 1 0 41124 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1649977179
transform 1 0 48024 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _231_
timestamp 1649977179
transform 1 0 64860 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _232_
timestamp 1649977179
transform 1 0 61272 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _233_
timestamp 1649977179
transform 1 0 62468 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1649977179
transform 1 0 82156 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _235_
timestamp 1649977179
transform 1 0 82708 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1649977179
transform 1 0 60628 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1649977179
transform 1 0 61824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _238_
timestamp 1649977179
transform 1 0 79120 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1649977179
transform 1 0 79120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1649977179
transform 1 0 82156 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _241_
timestamp 1649977179
transform 1 0 82708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _242_
timestamp 1649977179
transform 1 0 65872 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _243_
timestamp 1649977179
transform 1 0 90068 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1649977179
transform 1 0 92184 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _245_
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _246_
timestamp 1649977179
transform 1 0 46000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _247_
timestamp 1649977179
transform 1 0 46276 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _248_
timestamp 1649977179
transform 1 0 45356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _249_
timestamp 1649977179
transform 1 0 49864 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _251_
timestamp 1649977179
transform 1 0 89884 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _252_
timestamp 1649977179
transform 1 0 91724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _253_
timestamp 1649977179
transform 1 0 64584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _254_
timestamp 1649977179
transform 1 0 58788 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _255_
timestamp 1649977179
transform 1 0 58328 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _256_
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1649977179
transform 1 0 32660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _258_
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1649977179
transform 1 0 32660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _260_
timestamp 1649977179
transform 1 0 71852 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1649977179
transform 1 0 73324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1649977179
transform 1 0 71852 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _263_
timestamp 1649977179
transform 1 0 73324 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  _264_
timestamp 1649977179
transform 1 0 63940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _265_
timestamp 1649977179
transform 1 0 94392 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 1649977179
transform 1 0 95588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _267_
timestamp 1649977179
transform 1 0 59892 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _268_
timestamp 1649977179
transform 1 0 60536 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _269_
timestamp 1649977179
transform 1 0 71576 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _270_
timestamp 1649977179
transform 1 0 71116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _271_
timestamp 1649977179
transform 1 0 94300 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _272_
timestamp 1649977179
transform 1 0 94300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _273_
timestamp 1649977179
transform 1 0 60628 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1649977179
transform 1 0 58788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp 1649977179
transform 1 0 31188 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _277_
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _278_
timestamp 1649977179
transform 1 0 6624 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _279_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _280_
timestamp 1649977179
transform 1 0 57776 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _281_
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _282_
timestamp 1649977179
transform 1 0 57040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _283_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 68632 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _284_
timestamp 1649977179
transform 1 0 66976 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _285_ ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 66792 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _286_
timestamp 1649977179
transform 1 0 68632 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _287_
timestamp 1649977179
transform 1 0 66240 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _288_
timestamp 1649977179
transform 1 0 66240 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _298_
timestamp 1649977179
transform 1 0 19780 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _299_
timestamp 1649977179
transform 1 0 60720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1649977179
transform 1 0 47472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _301_
timestamp 1649977179
transform 1 0 51336 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _302_
timestamp 1649977179
transform 1 0 74428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _303_
timestamp 1649977179
transform 1 0 64308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _304_
timestamp 1649977179
transform 1 0 107364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _305_
timestamp 1649977179
transform 1 0 92644 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _306_
timestamp 1649977179
transform 1 0 104604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1649977179
transform 1 0 72864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _308_
timestamp 1649977179
transform 1 0 101200 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1649977179
transform 1 0 79028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _310_
timestamp 1649977179
transform 1 0 45908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _312_
timestamp 1649977179
transform 1 0 7912 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _313_
timestamp 1649977179
transform 1 0 32476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _314_
timestamp 1649977179
transform 1 0 107088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1649977179
transform 1 0 35236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _317_
timestamp 1649977179
transform 1 0 91264 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1649977179
transform 1 0 10488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _319_
timestamp 1649977179
transform 1 0 113528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _320_
timestamp 1649977179
transform 1 0 70012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _321_
timestamp 1649977179
transform 1 0 83996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1649977179
transform 1 0 86756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _323_
timestamp 1649977179
transform 1 0 10120 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _324_
timestamp 1649977179
transform 1 0 9292 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _325_
timestamp 1649977179
transform 1 0 113528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _327_
timestamp 1649977179
transform 1 0 28704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _328_
timestamp 1649977179
transform 1 0 57868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1649977179
transform 1 0 20516 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _331_
timestamp 1649977179
transform 1 0 59432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1649977179
transform 1 0 47748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1649977179
transform 1 0 50324 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _334_
timestamp 1649977179
transform 1 0 75164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1649977179
transform 1 0 63848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1649977179
transform 1 0 106812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1649977179
transform 1 0 103500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _338_
timestamp 1649977179
transform 1 0 104604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _339_
timestamp 1649977179
transform 1 0 73692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1649977179
transform 1 0 117208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _341_
timestamp 1649977179
transform 1 0 79672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _342_
timestamp 1649977179
transform 1 0 46552 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1649977179
transform 1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1649977179
transform 1 0 108008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _347_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _348_
timestamp 1649977179
transform 1 0 34500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1649977179
transform 1 0 95496 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _350_
timestamp 1649977179
transform 1 0 30544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _351_
timestamp 1649977179
transform 1 0 114540 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _352_
timestamp 1649977179
transform 1 0 71116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1649977179
transform 1 0 85376 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _354_
timestamp 1649977179
transform 1 0 86112 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1649977179
transform 1 0 2668 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _357_
timestamp 1649977179
transform 1 0 114540 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _358_
timestamp 1649977179
transform 1 0 50600 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _359_
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _360_
timestamp 1649977179
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _361_
timestamp 1649977179
transform 1 0 29440 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1649977179
transform 1 0 70748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _363_
timestamp 1649977179
transform 1 0 66884 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  bus_arbiter_316 ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 117944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  bus_arbiter_317
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  bus_arbiter_318
timestamp 1649977179
transform 1 0 115368 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  bus_arbiter_319
timestamp 1649977179
transform 1 0 99084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  bus_arbiter_320
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  bus_arbiter_321
timestamp 1649977179
transform 1 0 113436 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  bus_arbiter_322
timestamp 1649977179
transform 1 0 52256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  bus_arbiter_323
timestamp 1649977179
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  bus_arbiter_324
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk ~/hellochip/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 68540 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1649977179
transform 1 0 65044 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1649977179
transform 1 0 67620 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 74796 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1649977179
transform 1 0 6348 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 38456 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 43884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1649977179
transform 1 0 11500 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 27876 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform 1 0 33304 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform 1 0 117300 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 46828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 66884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 86204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1649977179
transform 1 0 117300 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1649977179
transform 1 0 81052 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 65044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 102488 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 59616 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1649977179
transform 1 0 116012 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1649977179
transform 1 0 111504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1649977179
transform 1 0 112148 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 77740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform 1 0 116288 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1649977179
transform 1 0 117668 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform 1 0 2392 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1649977179
transform 1 0 117300 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 72956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 66332 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 69092 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform 1 0 37628 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 68356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform 1 0 46736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1649977179
transform 1 0 28704 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1649977179
transform 1 0 100556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform 1 0 53544 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1649977179
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 40664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform 1 0 4968 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1649977179
transform 1 0 83628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform 1 0 59340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1649977179
transform 1 0 15548 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1649977179
transform 1 0 109756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 69644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform 1 0 79856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform 1 0 27140 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform 1 0 71852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform 1 0 86664 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1649977179
transform 1 0 82340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1649977179
transform 1 0 63204 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform 1 0 91540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1649977179
transform 1 0 15272 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform 1 0 77648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1649977179
transform 1 0 107180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1649977179
transform 1 0 117852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1649977179
transform 1 0 56488 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1649977179
transform 1 0 117852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform 1 0 117208 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1649977179
transform 1 0 105064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1649977179
transform 1 0 117116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1649977179
transform 1 0 49036 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1649977179
transform 1 0 117852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1649977179
transform 1 0 65596 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1649977179
transform 1 0 41676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1649977179
transform 1 0 61916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1649977179
transform 1 0 31280 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1649977179
transform 1 0 96876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1649977179
transform 1 0 12328 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input84
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1649977179
transform 1 0 36156 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1649977179
transform 1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1649977179
transform 1 0 117852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1649977179
transform 1 0 83628 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input90
timestamp 1649977179
transform 1 0 117484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input91
timestamp 1649977179
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input92
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1649977179
transform 1 0 116932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1649977179
transform 1 0 32476 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1649977179
transform 1 0 66240 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1649977179
transform 1 0 88780 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1649977179
transform 1 0 51980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input98
timestamp 1649977179
transform 1 0 117852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1649977179
transform 1 0 60812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1649977179
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input102
timestamp 1649977179
transform 1 0 91724 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1649977179
transform 1 0 117852 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1649977179
transform 1 0 97980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1649977179
transform 1 0 76084 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1649977179
transform 1 0 117116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1649977179
transform 1 0 117852 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input110
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1649977179
transform 1 0 89424 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1649977179
transform 1 0 75900 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input113
timestamp 1649977179
transform 1 0 7820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input114
timestamp 1649977179
transform 1 0 117668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input115
timestamp 1649977179
transform 1 0 76728 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input116
timestamp 1649977179
transform 1 0 87400 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input117
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input118
timestamp 1649977179
transform 1 0 102028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input119
timestamp 1649977179
transform 1 0 14260 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1649977179
transform 1 0 45816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1649977179
transform 1 0 112332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1649977179
transform 1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1649977179
transform 1 0 52900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input124
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input125
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input126
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1649977179
transform 1 0 101660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1649977179
transform 1 0 92184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1649977179
transform 1 0 21988 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input130
timestamp 1649977179
transform 1 0 99084 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input131
timestamp 1649977179
transform 1 0 117852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input133
timestamp 1649977179
transform 1 0 48024 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1649977179
transform 1 0 54556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input135
timestamp 1649977179
transform 1 0 17848 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input136
timestamp 1649977179
transform 1 0 25208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input137
timestamp 1649977179
transform 1 0 4140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input138
timestamp 1649977179
transform 1 0 72036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1649977179
transform 1 0 110860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1649977179
transform 1 0 61824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input141
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input142
timestamp 1649977179
transform 1 0 7544 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input143
timestamp 1649977179
transform 1 0 99452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input144
timestamp 1649977179
transform 1 0 81052 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input145
timestamp 1649977179
transform 1 0 117300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input146
timestamp 1649977179
transform 1 0 42412 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input147
timestamp 1649977179
transform 1 0 46460 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input150
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1649977179
transform 1 0 108100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input152
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1649977179
transform 1 0 105340 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input154
timestamp 1649977179
transform 1 0 117300 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input155
timestamp 1649977179
transform 1 0 59984 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input156
timestamp 1649977179
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input157
timestamp 1649977179
transform 1 0 114540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input158
timestamp 1649977179
transform 1 0 117852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input159
timestamp 1649977179
transform 1 0 26956 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input160
timestamp 1649977179
transform 1 0 117852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input161
timestamp 1649977179
transform 1 0 94760 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input162
timestamp 1649977179
transform 1 0 2668 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1649977179
transform 1 0 114540 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input164
timestamp 1649977179
transform 1 0 71944 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input165
timestamp 1649977179
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input166
timestamp 1649977179
transform 1 0 115368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input167
timestamp 1649977179
transform 1 0 58052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input168
timestamp 1649977179
transform 1 0 92828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input169
timestamp 1649977179
transform 1 0 20056 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input170
timestamp 1649977179
transform 1 0 74796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input171
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input172
timestamp 1649977179
transform 1 0 35512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input173
timestamp 1649977179
transform 1 0 103132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1649977179
transform 1 0 110032 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input175
timestamp 1649977179
transform 1 0 117852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input176
timestamp 1649977179
transform 1 0 110860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output177
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output178
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output179
timestamp 1649977179
transform 1 0 66792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output180
timestamp 1649977179
transform 1 0 79304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output181
timestamp 1649977179
transform 1 0 7820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output182
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output183
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output184
timestamp 1649977179
transform 1 0 105340 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output185
timestamp 1649977179
transform 1 0 81788 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output186
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output187
timestamp 1649977179
transform 1 0 36432 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output188
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output189
timestamp 1649977179
transform 1 0 105800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output190
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output191
timestamp 1649977179
transform 1 0 109388 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output192
timestamp 1649977179
transform 1 0 45816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output193
timestamp 1649977179
transform 1 0 84364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output194
timestamp 1649977179
transform 1 0 87032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output195
timestamp 1649977179
transform 1 0 10580 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output196
timestamp 1649977179
transform 1 0 93472 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output197
timestamp 1649977179
transform 1 0 102488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output198
timestamp 1649977179
transform 1 0 38088 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output199
timestamp 1649977179
transform 1 0 82524 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output200
timestamp 1649977179
transform 1 0 33580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output201
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output202
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output203
timestamp 1649977179
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output204
timestamp 1649977179
transform 1 0 38456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output205
timestamp 1649977179
transform 1 0 69368 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output206
timestamp 1649977179
transform 1 0 117944 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output207
timestamp 1649977179
transform 1 0 52900 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output208
timestamp 1649977179
transform 1 0 104420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output209
timestamp 1649977179
transform 1 0 73968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output210
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output211
timestamp 1649977179
transform 1 0 20792 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output212
timestamp 1649977179
transform 1 0 116380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output213
timestamp 1649977179
transform 1 0 117944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output214
timestamp 1649977179
transform 1 0 116012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output215
timestamp 1649977179
transform 1 0 56120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output216
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output217
timestamp 1649977179
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output218
timestamp 1649977179
transform 1 0 117944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output219
timestamp 1649977179
transform 1 0 97980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output220
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output221
timestamp 1649977179
transform 1 0 92828 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output222
timestamp 1649977179
transform 1 0 33396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output223
timestamp 1649977179
transform 1 0 56488 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output224
timestamp 1649977179
transform 1 0 117944 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output225
timestamp 1649977179
transform 1 0 71392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output226
timestamp 1649977179
transform 1 0 100556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output227
timestamp 1649977179
transform 1 0 4600 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output228
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output229
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output230
timestamp 1649977179
transform 1 0 117944 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output231
timestamp 1649977179
transform 1 0 50968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output232
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output233
timestamp 1649977179
transform 1 0 48392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output234
timestamp 1649977179
transform 1 0 95772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output235
timestamp 1649977179
transform 1 0 29716 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output236
timestamp 1649977179
transform 1 0 50968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output237
timestamp 1649977179
transform 1 0 95036 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output238
timestamp 1649977179
transform 1 0 64492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output239
timestamp 1649977179
transform 1 0 107456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output240
timestamp 1649977179
transform 1 0 116288 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output241
timestamp 1649977179
transform 1 0 77372 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output242
timestamp 1649977179
transform 1 0 50140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output243
timestamp 1649977179
transform 1 0 64492 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output244
timestamp 1649977179
transform 1 0 58696 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output245
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output246
timestamp 1649977179
transform 1 0 63204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output247
timestamp 1649977179
transform 1 0 87676 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output248
timestamp 1649977179
transform 1 0 117944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output249
timestamp 1649977179
transform 1 0 61824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output250
timestamp 1649977179
transform 1 0 84732 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output251
timestamp 1649977179
transform 1 0 90252 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output252
timestamp 1649977179
transform 1 0 78660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output253
timestamp 1649977179
transform 1 0 79764 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output254
timestamp 1649977179
transform 1 0 90252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output255
timestamp 1649977179
transform 1 0 111504 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output256
timestamp 1649977179
transform 1 0 97152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output257
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output258
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output259
timestamp 1649977179
transform 1 0 49956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output260
timestamp 1649977179
transform 1 0 117208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output261
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output262
timestamp 1649977179
transform 1 0 42596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output263
timestamp 1649977179
transform 1 0 46828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output264
timestamp 1649977179
transform 1 0 89608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output265
timestamp 1649977179
transform 1 0 65780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output266
timestamp 1649977179
transform 1 0 108284 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output267
timestamp 1649977179
transform 1 0 117944 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output268
timestamp 1649977179
transform 1 0 39376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output269
timestamp 1649977179
transform 1 0 55476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output270
timestamp 1649977179
transform 1 0 85100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output271
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output272
timestamp 1649977179
transform 1 0 37444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output273
timestamp 1649977179
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output274
timestamp 1649977179
transform 1 0 86204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output275
timestamp 1649977179
transform 1 0 110124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output276
timestamp 1649977179
transform 1 0 70748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output277
timestamp 1649977179
transform 1 0 88780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output278
timestamp 1649977179
transform 1 0 75900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output279
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output280
timestamp 1649977179
transform 1 0 113436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output281
timestamp 1649977179
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output282
timestamp 1649977179
transform 1 0 117944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output283
timestamp 1649977179
transform 1 0 106076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output284
timestamp 1649977179
transform 1 0 81236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output285
timestamp 1649977179
transform 1 0 103132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output286
timestamp 1649977179
transform 1 0 2668 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output287
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output288
timestamp 1649977179
transform 1 0 49036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output289
timestamp 1649977179
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output290
timestamp 1649977179
transform 1 0 57408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output291
timestamp 1649977179
transform 1 0 11684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output292
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output293
timestamp 1649977179
transform 1 0 70012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output294
timestamp 1649977179
transform 1 0 3312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output295
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output296
timestamp 1649977179
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output297
timestamp 1649977179
transform 1 0 87032 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output298
timestamp 1649977179
transform 1 0 70012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output299
timestamp 1649977179
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output300
timestamp 1649977179
transform 1 0 100372 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output301
timestamp 1649977179
transform 1 0 94116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output302
timestamp 1649977179
transform 1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output303
timestamp 1649977179
transform 1 0 117944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output304
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output305
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output306
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output307
timestamp 1649977179
transform 1 0 117944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output308
timestamp 1649977179
transform 1 0 44252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output309
timestamp 1649977179
transform 1 0 96508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output310
timestamp 1649977179
transform 1 0 95680 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output311
timestamp 1649977179
transform 1 0 41308 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output312
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output313
timestamp 1649977179
transform 1 0 53912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output314
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output315
timestamp 1649977179
transform 1 0 32936 0 -1 27200
box -38 -48 314 592
<< labels >>
flabel metal3 s 119200 8848 120000 8968 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 18694 29200 18750 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_ack_o
port 1 nsew signal tristate
flabel metal2 s 74722 29200 74778 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[0]
port 2 nsew signal input
flabel metal2 s 6458 29200 6514 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[10]
port 3 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[11]
port 4 nsew signal input
flabel metal2 s 39302 29200 39358 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[12]
port 5 nsew signal input
flabel metal2 s 43810 29200 43866 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[13]
port 6 nsew signal input
flabel metal2 s 10966 29200 11022 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[14]
port 7 nsew signal input
flabel metal2 s 28354 29200 28410 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[15]
port 8 nsew signal input
flabel metal2 s 33506 29200 33562 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[16]
port 9 nsew signal input
flabel metal3 s 119200 16328 120000 16448 0 FreeSans 480 0 0 0 m2_dcache_wbd_adr_i[17]
port 10 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[18]
port 11 nsew signal input
flabel metal2 s 66350 29200 66406 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[19]
port 12 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[1]
port 13 nsew signal input
flabel metal2 s 85670 0 85726 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[20]
port 14 nsew signal input
flabel metal3 s 119200 23128 120000 23248 0 FreeSans 480 0 0 0 m2_dcache_wbd_adr_i[21]
port 15 nsew signal input
flabel metal2 s 80518 0 80574 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[22]
port 16 nsew signal input
flabel metal2 s 64418 0 64474 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[23]
port 17 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[24]
port 18 nsew signal input
flabel metal2 s 102414 29200 102470 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[25]
port 19 nsew signal input
flabel metal2 s 59266 29200 59322 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[26]
port 20 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 m2_dcache_wbd_adr_i[27]
port 21 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 m2_dcache_wbd_adr_i[28]
port 22 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 m2_dcache_wbd_adr_i[29]
port 23 nsew signal input
flabel metal2 s 115938 29200 115994 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[2]
port 24 nsew signal input
flabel metal2 s 111430 0 111486 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[30]
port 25 nsew signal input
flabel metal2 s 112074 0 112130 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[31]
port 26 nsew signal input
flabel metal2 s 76654 0 76710 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[3]
port 27 nsew signal input
flabel metal3 s 119200 2048 120000 2168 0 FreeSans 480 0 0 0 m2_dcache_wbd_adr_i[4]
port 28 nsew signal input
flabel metal2 s 34794 29200 34850 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[5]
port 29 nsew signal input
flabel metal2 s 23846 29200 23902 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[6]
port 30 nsew signal input
flabel metal3 s 119200 4088 120000 4208 0 FreeSans 480 0 0 0 m2_dcache_wbd_adr_i[7]
port 31 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[8]
port 32 nsew signal input
flabel metal2 s 2594 29200 2650 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_adr_i[9]
port 33 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_cyc_i
port 34 nsew signal input
flabel metal3 s 119200 21088 120000 21208 0 FreeSans 480 0 0 0 m2_dcache_wbd_dat_i[0]
port 35 nsew signal input
flabel metal2 s 72790 29200 72846 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[10]
port 36 nsew signal input
flabel metal2 s 65706 29200 65762 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[11]
port 37 nsew signal input
flabel metal2 s 68282 29200 68338 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[12]
port 38 nsew signal input
flabel metal2 s 37370 29200 37426 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[13]
port 39 nsew signal input
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[14]
port 40 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[15]
port 41 nsew signal input
flabel metal2 s 28998 29200 29054 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[16]
port 42 nsew signal input
flabel metal2 s 100482 0 100538 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[17]
port 43 nsew signal input
flabel metal2 s 53470 29200 53526 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[18]
port 44 nsew signal input
flabel metal2 s 9034 29200 9090 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[19]
port 45 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[1]
port 46 nsew signal input
flabel metal2 s 5170 29200 5226 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[20]
port 47 nsew signal input
flabel metal2 s 13542 29200 13598 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[21]
port 48 nsew signal input
flabel metal2 s 83094 0 83150 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[22]
port 49 nsew signal input
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[23]
port 50 nsew signal input
flabel metal2 s 74078 0 74134 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[24]
port 51 nsew signal input
flabel metal2 s 15474 29200 15530 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[25]
port 52 nsew signal input
flabel metal2 s 108854 0 108910 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[26]
port 53 nsew signal input
flabel metal2 s 69570 0 69626 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[27]
port 54 nsew signal input
flabel metal2 s 78586 29200 78642 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[28]
port 55 nsew signal input
flabel metal2 s 27066 29200 27122 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[29]
port 56 nsew signal input
flabel metal2 s 70858 29200 70914 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[2]
port 57 nsew signal input
flabel metal2 s 85670 29200 85726 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[30]
port 58 nsew signal input
flabel metal2 s 81806 0 81862 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[31]
port 59 nsew signal input
flabel metal2 s 63130 29200 63186 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[3]
port 60 nsew signal input
flabel metal2 s 91466 0 91522 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[4]
port 61 nsew signal input
flabel metal2 s 16118 29200 16174 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[5]
port 62 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 m2_dcache_wbd_dat_i[6]
port 63 nsew signal input
flabel metal2 s 77298 0 77354 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[7]
port 64 nsew signal input
flabel metal2 s 106922 29200 106978 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_i[8]
port 65 nsew signal input
flabel metal3 s 119200 2728 120000 2848 0 FreeSans 480 0 0 0 m2_dcache_wbd_dat_i[9]
port 66 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[0]
port 67 nsew signal tristate
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[10]
port 68 nsew signal tristate
flabel metal2 s 79230 0 79286 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[11]
port 69 nsew signal tristate
flabel metal2 s 7746 29200 7802 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[12]
port 70 nsew signal tristate
flabel metal2 s 57334 29200 57390 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[13]
port 71 nsew signal tristate
flabel metal2 s 42522 29200 42578 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[14]
port 72 nsew signal tristate
flabel metal2 s 104346 29200 104402 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[15]
port 73 nsew signal tristate
flabel metal2 s 81162 29200 81218 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[16]
port 74 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 m2_dcache_wbd_dat_o[17]
port 75 nsew signal tristate
flabel metal2 s 35438 29200 35494 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[18]
port 76 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[19]
port 77 nsew signal tristate
flabel metal2 s 105634 0 105690 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[1]
port 78 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 m2_dcache_wbd_dat_o[20]
port 79 nsew signal tristate
flabel metal2 s 108854 29200 108910 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[21]
port 80 nsew signal tristate
flabel metal2 s 45742 29200 45798 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[22]
port 81 nsew signal tristate
flabel metal2 s 83738 0 83794 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[23]
port 82 nsew signal tristate
flabel metal2 s 86958 0 87014 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[24]
port 83 nsew signal tristate
flabel metal2 s 9678 29200 9734 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[25]
port 84 nsew signal tristate
flabel metal2 s 93398 29200 93454 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[26]
port 85 nsew signal tristate
flabel metal2 s 102414 0 102470 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[27]
port 86 nsew signal tristate
flabel metal2 s 38014 29200 38070 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[28]
port 87 nsew signal tristate
flabel metal2 s 82450 29200 82506 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[29]
port 88 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[2]
port 89 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 m2_dcache_wbd_dat_o[30]
port 90 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[31]
port 91 nsew signal tristate
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[3]
port 92 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[4]
port 93 nsew signal tristate
flabel metal2 s 67638 29200 67694 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[5]
port 94 nsew signal tristate
flabel metal3 s 119200 25168 120000 25288 0 FreeSans 480 0 0 0 m2_dcache_wbd_dat_o[6]
port 95 nsew signal tristate
flabel metal2 s 52826 29200 52882 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[7]
port 96 nsew signal tristate
flabel metal2 s 104346 0 104402 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[8]
port 97 nsew signal tristate
flabel metal2 s 72790 0 72846 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_dat_o[9]
port 98 nsew signal tristate
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_sel_i[0]
port 99 nsew signal input
flabel metal2 s 119802 0 119858 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_sel_i[1]
port 100 nsew signal input
flabel metal2 s 117870 29200 117926 30000 0 FreeSans 224 90 0 0 m2_dcache_wbd_sel_i[2]
port 101 nsew signal input
flabel metal2 s 104990 0 105046 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_sel_i[3]
port 102 nsew signal input
flabel metal3 s 119200 27888 120000 28008 0 FreeSans 480 0 0 0 m2_dcache_wbd_stb_i
port 103 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 m2_dcache_wbd_we_i
port 104 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 m2_others_wbd_ack_o
port 105 nsew signal tristate
flabel metal2 s 48962 29200 49018 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[0]
port 106 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 m2_others_wbd_adr_i[10]
port 107 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 m2_others_wbd_adr_i[11]
port 108 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[12]
port 109 nsew signal input
flabel metal3 s 119200 14288 120000 14408 0 FreeSans 480 0 0 0 m2_others_wbd_adr_i[13]
port 110 nsew signal input
flabel metal2 s 63774 29200 63830 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[14]
port 111 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[15]
port 112 nsew signal input
flabel metal2 s 61842 0 61898 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[16]
port 113 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[17]
port 114 nsew signal input
flabel metal2 s 30930 29200 30986 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[18]
port 115 nsew signal input
flabel metal2 s 96618 0 96674 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[19]
port 116 nsew signal input
flabel metal2 s 12254 29200 12310 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[1]
port 117 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 m2_others_wbd_adr_i[20]
port 118 nsew signal input
flabel metal2 s 36082 29200 36138 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[21]
port 119 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[22]
port 120 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 m2_others_wbd_adr_i[23]
port 121 nsew signal input
flabel metal3 s 119200 6128 120000 6248 0 FreeSans 480 0 0 0 m2_others_wbd_adr_i[24]
port 122 nsew signal input
flabel metal2 s 83094 29200 83150 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[25]
port 123 nsew signal input
flabel metal2 s 116582 0 116638 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[26]
port 124 nsew signal input
flabel metal2 s 17406 29200 17462 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[27]
port 125 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 m2_others_wbd_adr_i[28]
port 126 nsew signal input
flabel metal2 s 118514 0 118570 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[29]
port 127 nsew signal input
flabel metal2 s 31574 29200 31630 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[2]
port 128 nsew signal input
flabel metal2 s 64418 29200 64474 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[30]
port 129 nsew signal input
flabel metal2 s 88246 29200 88302 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[31]
port 130 nsew signal input
flabel metal2 s 52182 29200 52238 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[3]
port 131 nsew signal input
flabel metal3 s 119200 13608 120000 13728 0 FreeSans 480 0 0 0 m2_others_wbd_adr_i[4]
port 132 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[5]
port 133 nsew signal input
flabel metal2 s 59910 0 59966 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[6]
port 134 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[7]
port 135 nsew signal input
flabel metal2 s 91466 29200 91522 30000 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[8]
port 136 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 m2_others_wbd_adr_i[9]
port 137 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 m2_others_wbd_cyc_i
port 138 nsew signal input
flabel metal2 s 118514 29200 118570 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[0]
port 139 nsew signal input
flabel metal2 s 97906 0 97962 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[10]
port 140 nsew signal input
flabel metal2 s 76010 29200 76066 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[11]
port 141 nsew signal input
flabel metal3 s 119200 29248 120000 29368 0 FreeSans 480 0 0 0 m2_others_wbd_dat_i[12]
port 142 nsew signal input
flabel metal2 s 119802 29200 119858 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[13]
port 143 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 m2_others_wbd_dat_i[14]
port 144 nsew signal input
flabel metal2 s 89534 29200 89590 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[15]
port 145 nsew signal input
flabel metal2 s 74078 29200 74134 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[16]
port 146 nsew signal input
flabel metal2 s 7102 29200 7158 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[17]
port 147 nsew signal input
flabel metal3 s 119200 8 120000 128 0 FreeSans 480 0 0 0 m2_others_wbd_dat_i[18]
port 148 nsew signal input
flabel metal2 s 76654 29200 76710 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[19]
port 149 nsew signal input
flabel metal2 s 87602 0 87658 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[1]
port 150 nsew signal input
flabel metal2 s 1306 29200 1362 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[20]
port 151 nsew signal input
flabel metal2 s 101126 0 101182 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[21]
port 152 nsew signal input
flabel metal2 s 14186 29200 14242 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[22]
port 153 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[23]
port 154 nsew signal input
flabel metal2 s 112074 29200 112130 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[24]
port 155 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[25]
port 156 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[26]
port 157 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[27]
port 158 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[28]
port 159 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 m2_others_wbd_dat_i[29]
port 160 nsew signal input
flabel metal2 s 101126 29200 101182 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[2]
port 161 nsew signal input
flabel metal2 s 92110 0 92166 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[30]
port 162 nsew signal input
flabel metal2 s 21914 29200 21970 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[31]
port 163 nsew signal input
flabel metal2 s 98550 29200 98606 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[3]
port 164 nsew signal input
flabel metal3 s 119200 18368 120000 18488 0 FreeSans 480 0 0 0 m2_others_wbd_dat_i[4]
port 165 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[5]
port 166 nsew signal input
flabel metal2 s 48318 29200 48374 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[6]
port 167 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[7]
port 168 nsew signal input
flabel metal2 s 18050 29200 18106 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[8]
port 169 nsew signal input
flabel metal2 s 25134 29200 25190 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_i[9]
port 170 nsew signal input
flabel metal2 s 20626 29200 20682 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[0]
port 171 nsew signal tristate
flabel metal3 s 119200 1368 120000 1488 0 FreeSans 480 0 0 0 m2_others_wbd_dat_o[10]
port 172 nsew signal tristate
flabel metal3 s 119200 4768 120000 4888 0 FreeSans 480 0 0 0 m2_others_wbd_dat_o[11]
port 173 nsew signal tristate
flabel metal2 s 115938 0 115994 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[12]
port 174 nsew signal tristate
flabel metal2 s 55402 29200 55458 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[13]
port 175 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 m2_others_wbd_dat_o[14]
port 176 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[15]
port 177 nsew signal tristate
flabel metal3 s 119200 12928 120000 13048 0 FreeSans 480 0 0 0 m2_others_wbd_dat_o[16]
port 178 nsew signal tristate
flabel metal2 s 97906 29200 97962 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[17]
port 179 nsew signal tristate
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 m2_others_wbd_dat_o[18]
port 180 nsew signal tristate
flabel metal2 s 92110 29200 92166 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[19]
port 181 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[1]
port 182 nsew signal tristate
flabel metal2 s 56690 29200 56746 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[20]
port 183 nsew signal tristate
flabel metal3 s 119200 9528 120000 9648 0 FreeSans 480 0 0 0 m2_others_wbd_dat_o[21]
port 184 nsew signal tristate
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[22]
port 185 nsew signal tristate
flabel metal2 s 100482 29200 100538 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[23]
port 186 nsew signal tristate
flabel metal2 s 4526 29200 4582 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[24]
port 187 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[25]
port 188 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 m2_others_wbd_dat_o[26]
port 189 nsew signal tristate
flabel metal3 s 119200 20408 120000 20528 0 FreeSans 480 0 0 0 m2_others_wbd_dat_o[27]
port 190 nsew signal tristate
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[28]
port 191 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[29]
port 192 nsew signal tristate
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[2]
port 193 nsew signal tristate
flabel metal2 s 95974 0 96030 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[30]
port 194 nsew signal tristate
flabel metal2 s 29642 29200 29698 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[31]
port 195 nsew signal tristate
flabel metal2 s 50894 29200 50950 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[3]
port 196 nsew signal tristate
flabel metal2 s 94042 29200 94098 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[4]
port 197 nsew signal tristate
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[5]
port 198 nsew signal tristate
flabel metal2 s 106922 0 106978 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[6]
port 199 nsew signal tristate
flabel metal2 s 117226 29200 117282 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[7]
port 200 nsew signal tristate
flabel metal2 s 77298 29200 77354 30000 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[8]
port 201 nsew signal tristate
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 m2_others_wbd_dat_o[9]
port 202 nsew signal tristate
flabel metal2 s 3238 29200 3294 30000 0 FreeSans 224 90 0 0 m2_others_wbd_sel_i[0]
port 203 nsew signal input
flabel metal2 s 72146 0 72202 800 0 FreeSans 224 90 0 0 m2_others_wbd_sel_i[1]
port 204 nsew signal input
flabel metal2 s 110786 29200 110842 30000 0 FreeSans 224 90 0 0 m2_others_wbd_sel_i[2]
port 205 nsew signal input
flabel metal2 s 61198 0 61254 800 0 FreeSans 224 90 0 0 m2_others_wbd_sel_i[3]
port 206 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 m2_others_wbd_stb_i
port 207 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 m2_others_wbd_we_i
port 208 nsew signal input
flabel metal2 s 99194 0 99250 800 0 FreeSans 224 90 0 0 m2_wbd_ack_i
port 209 nsew signal input
flabel metal2 s 61842 29200 61898 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[0]
port 210 nsew signal tristate
flabel metal2 s 58622 29200 58678 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[10]
port 211 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 m2_wbd_adr_o[11]
port 212 nsew signal tristate
flabel metal2 s 63130 0 63186 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[12]
port 213 nsew signal tristate
flabel metal2 s 87602 29200 87658 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[13]
port 214 nsew signal tristate
flabel metal3 s 119200 24488 120000 24608 0 FreeSans 480 0 0 0 m2_wbd_adr_o[14]
port 215 nsew signal tristate
flabel metal2 s 61198 29200 61254 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[15]
port 216 nsew signal tristate
flabel metal2 s 83738 29200 83794 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[16]
port 217 nsew signal tristate
flabel metal2 s 90178 29200 90234 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[17]
port 218 nsew signal tristate
flabel metal2 s 78586 0 78642 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[18]
port 219 nsew signal tristate
flabel metal2 s 79230 29200 79286 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[19]
port 220 nsew signal tristate
flabel metal2 s 90178 0 90234 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[1]
port 221 nsew signal tristate
flabel metal2 s 111430 29200 111486 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[20]
port 222 nsew signal tristate
flabel metal2 s 96618 29200 96674 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[21]
port 223 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 m2_wbd_adr_o[22]
port 224 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[23]
port 225 nsew signal tristate
flabel metal2 s 50250 29200 50306 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[24]
port 226 nsew signal tristate
flabel metal2 s 117870 0 117926 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[25]
port 227 nsew signal tristate
flabel metal2 s 24490 29200 24546 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[26]
port 228 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[27]
port 229 nsew signal tristate
flabel metal2 s 47030 29200 47086 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[28]
port 230 nsew signal tristate
flabel metal2 s 89534 0 89590 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[29]
port 231 nsew signal tristate
flabel metal2 s 65706 0 65762 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[2]
port 232 nsew signal tristate
flabel metal2 s 107566 29200 107622 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[30]
port 233 nsew signal tristate
flabel metal3 s 119200 22448 120000 22568 0 FreeSans 480 0 0 0 m2_wbd_adr_o[31]
port 234 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[3]
port 235 nsew signal tristate
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[4]
port 236 nsew signal tristate
flabel metal2 s 85026 0 85082 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[5]
port 237 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 m2_wbd_adr_o[6]
port 238 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[7]
port 239 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 m2_wbd_adr_o[8]
port 240 nsew signal tristate
flabel metal2 s 85026 29200 85082 30000 0 FreeSans 224 90 0 0 m2_wbd_adr_o[9]
port 241 nsew signal tristate
flabel metal2 s 109498 0 109554 800 0 FreeSans 224 90 0 0 m2_wbd_bl_o[0]
port 242 nsew signal tristate
flabel metal3 s 119200 15648 120000 15768 0 FreeSans 480 0 0 0 m2_wbd_bl_o[1]
port 243 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 m2_wbd_bl_o[2]
port 244 nsew signal tristate
flabel metal2 s 115294 29200 115350 30000 0 FreeSans 224 90 0 0 m2_wbd_bl_o[3]
port 245 nsew signal tristate
flabel metal2 s 98550 0 98606 800 0 FreeSans 224 90 0 0 m2_wbd_bl_o[4]
port 246 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 m2_wbd_bl_o[5]
port 247 nsew signal tristate
flabel metal2 s 113362 29200 113418 30000 0 FreeSans 224 90 0 0 m2_wbd_bl_o[6]
port 248 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 m2_wbd_bl_o[7]
port 249 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 m2_wbd_bl_o[8]
port 250 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 m2_wbd_bl_o[9]
port 251 nsew signal tristate
flabel metal2 s 70214 0 70270 800 0 FreeSans 224 90 0 0 m2_wbd_bry_o
port 252 nsew signal tristate
flabel metal2 s 88246 0 88302 800 0 FreeSans 224 90 0 0 m2_wbd_cyc_o
port 253 nsew signal tristate
flabel metal2 s 80518 29200 80574 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[0]
port 254 nsew signal input
flabel metal3 s 119200 11568 120000 11688 0 FreeSans 480 0 0 0 m2_wbd_dat_i[10]
port 255 nsew signal input
flabel metal2 s 41878 29200 41934 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[11]
port 256 nsew signal input
flabel metal2 s 46386 29200 46442 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[12]
port 257 nsew signal input
flabel metal2 s 44454 29200 44510 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[13]
port 258 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[14]
port 259 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[15]
port 260 nsew signal input
flabel metal2 s 107566 0 107622 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[16]
port 261 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 m2_wbd_dat_i[17]
port 262 nsew signal input
flabel metal2 s 104990 29200 105046 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[18]
port 263 nsew signal input
flabel metal3 s 119200 27208 120000 27328 0 FreeSans 480 0 0 0 m2_wbd_dat_i[19]
port 264 nsew signal input
flabel metal2 s 59910 29200 59966 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[1]
port 265 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[20]
port 266 nsew signal input
flabel metal2 s 114006 0 114062 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[21]
port 267 nsew signal input
flabel metal3 s 119200 26528 120000 26648 0 FreeSans 480 0 0 0 m2_wbd_dat_i[22]
port 268 nsew signal input
flabel metal2 s 26422 29200 26478 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[23]
port 269 nsew signal input
flabel metal3 s 119200 6808 120000 6928 0 FreeSans 480 0 0 0 m2_wbd_dat_i[24]
port 270 nsew signal input
flabel metal2 s 94686 0 94742 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[25]
port 271 nsew signal input
flabel metal2 s 18 29200 74 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[26]
port 272 nsew signal input
flabel metal2 s 114006 29200 114062 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[27]
port 273 nsew signal input
flabel metal2 s 72146 29200 72202 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[28]
port 274 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[29]
port 275 nsew signal input
flabel metal2 s 115294 0 115350 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[2]
port 276 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[30]
port 277 nsew signal input
flabel metal2 s 92754 0 92810 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[31]
port 278 nsew signal input
flabel metal2 s 19982 29200 20038 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[3]
port 279 nsew signal input
flabel metal2 s 74722 0 74778 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[4]
port 280 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[5]
port 281 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[6]
port 282 nsew signal input
flabel metal2 s 103058 0 103114 800 0 FreeSans 224 90 0 0 m2_wbd_dat_i[7]
port 283 nsew signal input
flabel metal2 s 109498 29200 109554 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_i[8]
port 284 nsew signal input
flabel metal3 s 119200 17688 120000 17808 0 FreeSans 480 0 0 0 m2_wbd_dat_i[9]
port 285 nsew signal input
flabel metal2 s 75366 0 75422 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[0]
port 286 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 m2_wbd_dat_o[10]
port 287 nsew signal tristate
flabel metal2 s 113362 0 113418 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[11]
port 288 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[12]
port 289 nsew signal tristate
flabel metal3 s 119200 19728 120000 19848 0 FreeSans 480 0 0 0 m2_wbd_dat_o[13]
port 290 nsew signal tristate
flabel metal2 s 105634 29200 105690 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[14]
port 291 nsew signal tristate
flabel metal2 s 81162 0 81218 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[15]
port 292 nsew signal tristate
flabel metal2 s 103058 29200 103114 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[16]
port 293 nsew signal tristate
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 m2_wbd_dat_o[17]
port 294 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 m2_wbd_dat_o[18]
port 295 nsew signal tristate
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[19]
port 296 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[1]
port 297 nsew signal tristate
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[20]
port 298 nsew signal tristate
flabel metal2 s 11610 29200 11666 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[21]
port 299 nsew signal tristate
flabel metal2 s 39946 29200 40002 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[22]
port 300 nsew signal tristate
flabel metal2 s 69570 29200 69626 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[23]
port 301 nsew signal tristate
flabel metal2 s 662 29200 718 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[24]
port 302 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[25]
port 303 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[26]
port 304 nsew signal tristate
flabel metal2 s 86958 29200 87014 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[27]
port 305 nsew signal tristate
flabel metal2 s 70214 29200 70270 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[28]
port 306 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[29]
port 307 nsew signal tristate
flabel metal2 s 99838 29200 99894 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[2]
port 308 nsew signal tristate
flabel metal2 s 94042 0 94098 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[30]
port 309 nsew signal tristate
flabel metal2 s 22558 29200 22614 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[31]
port 310 nsew signal tristate
flabel metal3 s 119200 10888 120000 11008 0 FreeSans 480 0 0 0 m2_wbd_dat_o[3]
port 311 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[4]
port 312 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[5]
port 313 nsew signal tristate
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 m2_wbd_dat_o[6]
port 314 nsew signal tristate
flabel metal3 s 119200 8168 120000 8288 0 FreeSans 480 0 0 0 m2_wbd_dat_o[7]
port 315 nsew signal tristate
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 m2_wbd_dat_o[8]
port 316 nsew signal tristate
flabel metal2 s 95974 29200 96030 30000 0 FreeSans 224 90 0 0 m2_wbd_dat_o[9]
port 317 nsew signal tristate
flabel metal2 s 94686 29200 94742 30000 0 FreeSans 224 90 0 0 m2_wbd_sel_o[0]
port 318 nsew signal tristate
flabel metal2 s 41234 29200 41290 30000 0 FreeSans 224 90 0 0 m2_wbd_sel_o[1]
port 319 nsew signal tristate
flabel metal2 s 54758 29200 54814 30000 0 FreeSans 224 90 0 0 m2_wbd_sel_o[2]
port 320 nsew signal tristate
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 m2_wbd_sel_o[3]
port 321 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 m2_wbd_stb_o
port 322 nsew signal tristate
flabel metal2 s 32862 29200 32918 30000 0 FreeSans 224 90 0 0 m2_wbd_we_o
port 323 nsew signal tristate
flabel metal2 s 110786 0 110842 800 0 FreeSans 224 90 0 0 reset
port 324 nsew signal input
flabel metal4 s 15668 2128 15988 27792 0 FreeSans 1920 90 0 0 vccd1
port 325 nsew power bidirectional
flabel metal4 s 45116 2128 45436 27792 0 FreeSans 1920 90 0 0 vccd1
port 325 nsew power bidirectional
flabel metal4 s 74564 2128 74884 27792 0 FreeSans 1920 90 0 0 vccd1
port 325 nsew power bidirectional
flabel metal4 s 104012 2128 104332 27792 0 FreeSans 1920 90 0 0 vccd1
port 325 nsew power bidirectional
flabel metal4 s 30392 2128 30712 27792 0 FreeSans 1920 90 0 0 vssd1
port 326 nsew ground bidirectional
flabel metal4 s 59840 2128 60160 27792 0 FreeSans 1920 90 0 0 vssd1
port 326 nsew ground bidirectional
flabel metal4 s 89288 2128 89608 27792 0 FreeSans 1920 90 0 0 vssd1
port 326 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 30000
<< end >>
