VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO l1icache_32
  CLASS BLOCK ;
  FOREIGN l1icache_32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 150.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END clk
  PIN data_chip_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 146.000 26.130 150.000 ;
    END
  END data_chip_en
  PIN data_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 37.440 450.000 38.040 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 146.000 177.470 150.000 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 57.840 450.000 58.440 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 146.000 74.430 150.000 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 146.000 361.010 150.000 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 146.000 212.890 150.000 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 146.000 174.250 150.000 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 146.000 51.890 150.000 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 146.000 261.190 150.000 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 146.000 3.590 150.000 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 146.000 0.370 150.000 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 146.000 309.490 150.000 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 146.000 228.990 150.000 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 146.000 357.790 150.000 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 146.000 167.810 150.000 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 146.000 100.190 150.000 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END data_in[31]
  PIN data_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 146.000 325.590 150.000 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 146.000 35.790 150.000 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 146.000 193.570 150.000 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 146.000 196.790 150.000 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 146.000 386.770 150.000 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END data_in[9]
  PIN data_index[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 146.000 180.690 150.000 ;
    END
  END data_index[0]
  PIN data_index[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 105.440 450.000 106.040 ;
    END
  END data_index[1]
  PIN data_index[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 146.000 409.310 150.000 ;
    END
  END data_index[2]
  PIN data_index[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 142.840 450.000 143.440 ;
    END
  END data_index[3]
  PIN data_index[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END data_index[4]
  PIN data_index[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 146.000 77.650 150.000 ;
    END
  END data_index[5]
  PIN data_index[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 146.000 370.670 150.000 ;
    END
  END data_index[6]
  PIN data_index[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END data_index[7]
  PIN data_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 146.000 80.870 150.000 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 132.640 450.000 133.240 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 146.000 64.770 150.000 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 146.000 209.670 150.000 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 44.240 450.000 44.840 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 146.000 32.570 150.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 146.000 58.330 150.000 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 146.000 438.290 150.000 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 40.840 450.000 41.440 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 146.000 418.970 150.000 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 146.000 119.510 150.000 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 146.000 106.630 150.000 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 146.000 425.410 150.000 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 146.000 22.910 150.000 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 34.040 450.000 34.640 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 146.000 257.970 150.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 54.440 450.000 55.040 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 146.000 154.930 150.000 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 146.000 270.850 150.000 ;
    END
  END data_out[9]
  PIN data_write_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 146.000 441.510 150.000 ;
    END
  END data_write_en
  PIN ld_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END ld_data_o[0]
  PIN ld_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 146.000 373.890 150.000 ;
    END
  END ld_data_o[10]
  PIN ld_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 13.640 450.000 14.240 ;
    END
  END ld_data_o[11]
  PIN ld_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END ld_data_o[12]
  PIN ld_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 146.000 219.330 150.000 ;
    END
  END ld_data_o[13]
  PIN ld_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END ld_data_o[14]
  PIN ld_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 95.240 450.000 95.840 ;
    END
  END ld_data_o[15]
  PIN ld_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 146.000 225.770 150.000 ;
    END
  END ld_data_o[16]
  PIN ld_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END ld_data_o[17]
  PIN ld_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 146.000 45.450 150.000 ;
    END
  END ld_data_o[18]
  PIN ld_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END ld_data_o[19]
  PIN ld_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 68.040 450.000 68.640 ;
    END
  END ld_data_o[1]
  PIN ld_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 146.000 364.230 150.000 ;
    END
  END ld_data_o[20]
  PIN ld_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END ld_data_o[21]
  PIN ld_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 23.840 450.000 24.440 ;
    END
  END ld_data_o[22]
  PIN ld_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 146.000 444.730 150.000 ;
    END
  END ld_data_o[23]
  PIN ld_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 146.000 348.130 150.000 ;
    END
  END ld_data_o[24]
  PIN ld_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END ld_data_o[25]
  PIN ld_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 146.000 296.610 150.000 ;
    END
  END ld_data_o[26]
  PIN ld_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 20.440 450.000 21.040 ;
    END
  END ld_data_o[27]
  PIN ld_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END ld_data_o[28]
  PIN ld_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 146.000 435.070 150.000 ;
    END
  END ld_data_o[29]
  PIN ld_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 146.000 312.710 150.000 ;
    END
  END ld_data_o[2]
  PIN ld_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END ld_data_o[30]
  PIN ld_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END ld_data_o[31]
  PIN ld_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 0.040 450.000 0.640 ;
    END
  END ld_data_o[3]
  PIN ld_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END ld_data_o[4]
  PIN ld_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 146.000 254.750 150.000 ;
    END
  END ld_data_o[5]
  PIN ld_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END ld_data_o[6]
  PIN ld_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END ld_data_o[7]
  PIN ld_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END ld_data_o[8]
  PIN ld_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END ld_data_o[9]
  PIN req_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END req_addr_i[0]
  PIN req_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 146.000 399.650 150.000 ;
    END
  END req_addr_i[10]
  PIN req_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END req_addr_i[11]
  PIN req_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END req_addr_i[12]
  PIN req_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END req_addr_i[13]
  PIN req_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 146.000 222.550 150.000 ;
    END
  END req_addr_i[14]
  PIN req_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END req_addr_i[15]
  PIN req_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 146.000 145.270 150.000 ;
    END
  END req_addr_i[16]
  PIN req_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 146.000 113.070 150.000 ;
    END
  END req_addr_i[17]
  PIN req_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 146.000 335.250 150.000 ;
    END
  END req_addr_i[18]
  PIN req_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END req_addr_i[19]
  PIN req_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 146.000 267.630 150.000 ;
    END
  END req_addr_i[1]
  PIN req_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END req_addr_i[20]
  PIN req_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 30.640 450.000 31.240 ;
    END
  END req_addr_i[21]
  PIN req_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END req_addr_i[22]
  PIN req_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END req_addr_i[23]
  PIN req_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 91.840 450.000 92.440 ;
    END
  END req_addr_i[24]
  PIN req_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END req_addr_i[25]
  PIN req_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 146.000 183.910 150.000 ;
    END
  END req_addr_i[26]
  PIN req_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 146.000 142.050 150.000 ;
    END
  END req_addr_i[27]
  PIN req_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 146.000 84.090 150.000 ;
    END
  END req_addr_i[28]
  PIN req_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 146.000 412.530 150.000 ;
    END
  END req_addr_i[29]
  PIN req_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END req_addr_i[2]
  PIN req_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END req_addr_i[30]
  PIN req_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END req_addr_i[31]
  PIN req_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 146.000 6.810 150.000 ;
    END
  END req_addr_i[3]
  PIN req_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 146.000 447.950 150.000 ;
    END
  END req_addr_i[4]
  PIN req_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END req_addr_i[5]
  PIN req_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END req_addr_i[6]
  PIN req_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 146.000 116.290 150.000 ;
    END
  END req_addr_i[7]
  PIN req_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END req_addr_i[8]
  PIN req_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 146.000 338.470 150.000 ;
    END
  END req_addr_i[9]
  PIN req_ready_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 115.640 450.000 116.240 ;
    END
  END req_ready_o
  PIN req_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 146.000 341.690 150.000 ;
    END
  END req_valid_i
  PIN resp_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END resp_addr_o[0]
  PIN resp_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END resp_addr_o[10]
  PIN resp_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 146.000 109.850 150.000 ;
    END
  END resp_addr_o[11]
  PIN resp_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 108.840 450.000 109.440 ;
    END
  END resp_addr_o[12]
  PIN resp_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END resp_addr_o[13]
  PIN resp_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END resp_addr_o[14]
  PIN resp_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 146.000 377.110 150.000 ;
    END
  END resp_addr_o[15]
  PIN resp_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END resp_addr_o[16]
  PIN resp_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END resp_addr_o[17]
  PIN resp_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 146.000 283.730 150.000 ;
    END
  END resp_addr_o[18]
  PIN resp_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 146.000 428.630 150.000 ;
    END
  END resp_addr_o[19]
  PIN resp_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END resp_addr_o[1]
  PIN resp_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END resp_addr_o[20]
  PIN resp_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 146.000 245.090 150.000 ;
    END
  END resp_addr_o[21]
  PIN resp_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 81.640 450.000 82.240 ;
    END
  END resp_addr_o[22]
  PIN resp_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END resp_addr_o[23]
  PIN resp_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 146.000 328.810 150.000 ;
    END
  END resp_addr_o[24]
  PIN resp_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 146.000 303.050 150.000 ;
    END
  END resp_addr_o[25]
  PIN resp_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END resp_addr_o[26]
  PIN resp_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 146.000 280.510 150.000 ;
    END
  END resp_addr_o[27]
  PIN resp_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 146.000 206.450 150.000 ;
    END
  END resp_addr_o[28]
  PIN resp_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END resp_addr_o[29]
  PIN resp_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END resp_addr_o[2]
  PIN resp_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END resp_addr_o[30]
  PIN resp_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END resp_addr_o[31]
  PIN resp_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END resp_addr_o[3]
  PIN resp_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 146.000 232.210 150.000 ;
    END
  END resp_addr_o[4]
  PIN resp_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END resp_addr_o[5]
  PIN resp_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END resp_addr_o[6]
  PIN resp_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END resp_addr_o[7]
  PIN resp_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END resp_addr_o[8]
  PIN resp_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END resp_addr_o[9]
  PIN resp_ready_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END resp_ready_i
  PIN resp_valid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END resp_valid_o
  PIN rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 74.840 450.000 75.440 ;
    END
  END rstn
  PIN tag_chip_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 146.000 216.110 150.000 ;
    END
  END tag_chip_en
  PIN tag_data_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END tag_data_in[0]
  PIN tag_data_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END tag_data_in[10]
  PIN tag_data_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END tag_data_in[11]
  PIN tag_data_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 146.000 171.030 150.000 ;
    END
  END tag_data_in[12]
  PIN tag_data_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 146.000 71.210 150.000 ;
    END
  END tag_data_in[13]
  PIN tag_data_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 146.000 13.250 150.000 ;
    END
  END tag_data_in[14]
  PIN tag_data_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END tag_data_in[15]
  PIN tag_data_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 51.040 450.000 51.640 ;
    END
  END tag_data_in[16]
  PIN tag_data_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END tag_data_in[17]
  PIN tag_data_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 146.000 164.590 150.000 ;
    END
  END tag_data_in[18]
  PIN tag_data_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END tag_data_in[19]
  PIN tag_data_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 17.040 450.000 17.640 ;
    END
  END tag_data_in[1]
  PIN tag_data_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END tag_data_in[20]
  PIN tag_data_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 98.640 450.000 99.240 ;
    END
  END tag_data_in[21]
  PIN tag_data_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END tag_data_in[22]
  PIN tag_data_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END tag_data_in[23]
  PIN tag_data_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 146.000 322.370 150.000 ;
    END
  END tag_data_in[24]
  PIN tag_data_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END tag_data_in[25]
  PIN tag_data_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END tag_data_in[26]
  PIN tag_data_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 85.040 450.000 85.640 ;
    END
  END tag_data_in[27]
  PIN tag_data_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END tag_data_in[28]
  PIN tag_data_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END tag_data_in[29]
  PIN tag_data_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 146.000 90.530 150.000 ;
    END
  END tag_data_in[2]
  PIN tag_data_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END tag_data_in[30]
  PIN tag_data_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END tag_data_in[31]
  PIN tag_data_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 122.440 450.000 123.040 ;
    END
  END tag_data_in[3]
  PIN tag_data_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 146.000 122.730 150.000 ;
    END
  END tag_data_in[4]
  PIN tag_data_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END tag_data_in[5]
  PIN tag_data_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 146.000 19.690 150.000 ;
    END
  END tag_data_in[6]
  PIN tag_data_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END tag_data_in[7]
  PIN tag_data_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 146.000 190.350 150.000 ;
    END
  END tag_data_in[8]
  PIN tag_data_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 146.000 290.170 150.000 ;
    END
  END tag_data_in[9]
  PIN tag_index[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 146.000 332.030 150.000 ;
    END
  END tag_index[0]
  PIN tag_index[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END tag_index[1]
  PIN tag_index[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END tag_index[2]
  PIN tag_index[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 146.000 93.750 150.000 ;
    END
  END tag_index[3]
  PIN tag_index[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 146.000 264.410 150.000 ;
    END
  END tag_index[4]
  PIN tag_index[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END tag_index[5]
  PIN tag_index[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 119.040 450.000 119.640 ;
    END
  END tag_index[6]
  PIN tag_index[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END tag_index[7]
  PIN tag_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 146.000 396.430 150.000 ;
    END
  END tag_out[0]
  PIN tag_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END tag_out[10]
  PIN tag_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 146.000 151.710 150.000 ;
    END
  END tag_out[11]
  PIN tag_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END tag_out[12]
  PIN tag_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END tag_out[13]
  PIN tag_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 146.000 158.150 150.000 ;
    END
  END tag_out[14]
  PIN tag_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END tag_out[15]
  PIN tag_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END tag_out[16]
  PIN tag_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END tag_out[17]
  PIN tag_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 146.000 306.270 150.000 ;
    END
  END tag_out[18]
  PIN tag_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 136.040 450.000 136.640 ;
    END
  END tag_out[19]
  PIN tag_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 146.000 55.110 150.000 ;
    END
  END tag_out[1]
  PIN tag_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 146.000 293.390 150.000 ;
    END
  END tag_out[20]
  PIN tag_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END tag_out[21]
  PIN tag_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END tag_out[22]
  PIN tag_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 146.000 274.070 150.000 ;
    END
  END tag_out[23]
  PIN tag_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END tag_out[24]
  PIN tag_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 146.000 402.870 150.000 ;
    END
  END tag_out[25]
  PIN tag_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END tag_out[26]
  PIN tag_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 146.000 235.430 150.000 ;
    END
  END tag_out[27]
  PIN tag_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END tag_out[28]
  PIN tag_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END tag_out[29]
  PIN tag_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 27.240 450.000 27.840 ;
    END
  END tag_out[2]
  PIN tag_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 146.000 29.350 150.000 ;
    END
  END tag_out[30]
  PIN tag_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END tag_out[31]
  PIN tag_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 146.000 96.970 150.000 ;
    END
  END tag_out[3]
  PIN tag_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END tag_out[4]
  PIN tag_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END tag_out[5]
  PIN tag_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END tag_out[6]
  PIN tag_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 125.840 450.000 126.440 ;
    END
  END tag_out[7]
  PIN tag_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END tag_out[8]
  PIN tag_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END tag_out[9]
  PIN tag_write_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END tag_write_en
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 59.590 10.640 61.190 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.330 10.640 170.930 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.070 10.640 280.670 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 388.810 10.640 390.410 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 114.460 10.640 116.060 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.200 10.640 225.800 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 333.940 10.640 335.540 138.960 ;
    END
  END vssd1
  PIN wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 146.000 241.870 150.000 ;
    END
  END wb_ack_i
  PIN wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wb_adr_o[0]
  PIN wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wb_adr_o[10]
  PIN wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 146.000 299.830 150.000 ;
    END
  END wb_adr_o[11]
  PIN wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END wb_adr_o[12]
  PIN wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END wb_adr_o[13]
  PIN wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wb_adr_o[14]
  PIN wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 146.000 39.010 150.000 ;
    END
  END wb_adr_o[15]
  PIN wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END wb_adr_o[16]
  PIN wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END wb_adr_o[17]
  PIN wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 146.000 415.750 150.000 ;
    END
  END wb_adr_o[18]
  PIN wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END wb_adr_o[19]
  PIN wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wb_adr_o[1]
  PIN wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wb_adr_o[20]
  PIN wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END wb_adr_o[21]
  PIN wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END wb_adr_o[22]
  PIN wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 146.000 286.950 150.000 ;
    END
  END wb_adr_o[23]
  PIN wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 78.240 450.000 78.840 ;
    END
  END wb_adr_o[24]
  PIN wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 146.000 132.390 150.000 ;
    END
  END wb_adr_o[25]
  PIN wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 146.000 148.490 150.000 ;
    END
  END wb_adr_o[26]
  PIN wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 146.000 138.830 150.000 ;
    END
  END wb_adr_o[27]
  PIN wb_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END wb_adr_o[28]
  PIN wb_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wb_adr_o[29]
  PIN wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END wb_adr_o[2]
  PIN wb_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END wb_adr_o[30]
  PIN wb_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 146.000 383.550 150.000 ;
    END
  END wb_adr_o[31]
  PIN wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 146.240 450.000 146.840 ;
    END
  END wb_adr_o[3]
  PIN wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 146.000 203.230 150.000 ;
    END
  END wb_adr_o[4]
  PIN wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wb_adr_o[5]
  PIN wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wb_adr_o[6]
  PIN wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 139.440 450.000 140.040 ;
    END
  END wb_adr_o[7]
  PIN wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 146.000 67.990 150.000 ;
    END
  END wb_adr_o[8]
  PIN wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 61.240 450.000 61.840 ;
    END
  END wb_adr_o[9]
  PIN wb_bl_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END wb_bl_o[0]
  PIN wb_bl_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END wb_bl_o[1]
  PIN wb_bl_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 146.000 422.190 150.000 ;
    END
  END wb_bl_o[2]
  PIN wb_bl_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END wb_bl_o[3]
  PIN wb_bl_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wb_bl_o[4]
  PIN wb_bl_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 10.240 450.000 10.840 ;
    END
  END wb_bl_o[5]
  PIN wb_bl_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END wb_bl_o[6]
  PIN wb_bl_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END wb_bl_o[7]
  PIN wb_bl_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 146.000 42.230 150.000 ;
    END
  END wb_bl_o[8]
  PIN wb_bl_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wb_bl_o[9]
  PIN wb_bry_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wb_bry_o
  PIN wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wb_cyc_o
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 146.000 406.090 150.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 102.040 450.000 102.640 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 3.440 450.000 4.040 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 112.240 450.000 112.840 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 146.000 389.990 150.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 146.000 380.330 150.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 146.000 16.470 150.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 146.000 129.170 150.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 146.000 248.310 150.000 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 146.000 319.150 150.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 146.000 251.530 150.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 146.000 367.450 150.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 146.000 61.550 150.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 71.440 450.000 72.040 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wb_dat_i[9]
  PIN wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 64.640 450.000 65.240 ;
    END
  END wb_stb_o
  PIN wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wb_we_o
  PIN write_data_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 146.000 351.350 150.000 ;
    END
  END write_data_mask[0]
  PIN write_data_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 146.000 344.910 150.000 ;
    END
  END write_data_mask[1]
  PIN write_data_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 146.000 135.610 150.000 ;
    END
  END write_data_mask[2]
  PIN write_data_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 146.000 187.130 150.000 ;
    END
  END write_data_mask[3]
  PIN write_tag_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END write_tag_mask[0]
  PIN write_tag_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END write_tag_mask[1]
  PIN write_tag_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 146.000 103.410 150.000 ;
    END
  END write_tag_mask[2]
  PIN write_tag_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END write_tag_mask[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 444.360 138.805 ;
      LAYER met1 ;
        RECT 0.070 5.820 447.970 138.960 ;
      LAYER met2 ;
        RECT 0.650 145.720 3.030 146.725 ;
        RECT 3.870 145.720 6.250 146.725 ;
        RECT 7.090 145.720 12.690 146.725 ;
        RECT 13.530 145.720 15.910 146.725 ;
        RECT 16.750 145.720 19.130 146.725 ;
        RECT 19.970 145.720 22.350 146.725 ;
        RECT 23.190 145.720 25.570 146.725 ;
        RECT 26.410 145.720 28.790 146.725 ;
        RECT 29.630 145.720 32.010 146.725 ;
        RECT 32.850 145.720 35.230 146.725 ;
        RECT 36.070 145.720 38.450 146.725 ;
        RECT 39.290 145.720 41.670 146.725 ;
        RECT 42.510 145.720 44.890 146.725 ;
        RECT 45.730 145.720 51.330 146.725 ;
        RECT 52.170 145.720 54.550 146.725 ;
        RECT 55.390 145.720 57.770 146.725 ;
        RECT 58.610 145.720 60.990 146.725 ;
        RECT 61.830 145.720 64.210 146.725 ;
        RECT 65.050 145.720 67.430 146.725 ;
        RECT 68.270 145.720 70.650 146.725 ;
        RECT 71.490 145.720 73.870 146.725 ;
        RECT 74.710 145.720 77.090 146.725 ;
        RECT 77.930 145.720 80.310 146.725 ;
        RECT 81.150 145.720 83.530 146.725 ;
        RECT 84.370 145.720 89.970 146.725 ;
        RECT 90.810 145.720 93.190 146.725 ;
        RECT 94.030 145.720 96.410 146.725 ;
        RECT 97.250 145.720 99.630 146.725 ;
        RECT 100.470 145.720 102.850 146.725 ;
        RECT 103.690 145.720 106.070 146.725 ;
        RECT 106.910 145.720 109.290 146.725 ;
        RECT 110.130 145.720 112.510 146.725 ;
        RECT 113.350 145.720 115.730 146.725 ;
        RECT 116.570 145.720 118.950 146.725 ;
        RECT 119.790 145.720 122.170 146.725 ;
        RECT 123.010 145.720 128.610 146.725 ;
        RECT 129.450 145.720 131.830 146.725 ;
        RECT 132.670 145.720 135.050 146.725 ;
        RECT 135.890 145.720 138.270 146.725 ;
        RECT 139.110 145.720 141.490 146.725 ;
        RECT 142.330 145.720 144.710 146.725 ;
        RECT 145.550 145.720 147.930 146.725 ;
        RECT 148.770 145.720 151.150 146.725 ;
        RECT 151.990 145.720 154.370 146.725 ;
        RECT 155.210 145.720 157.590 146.725 ;
        RECT 158.430 145.720 164.030 146.725 ;
        RECT 164.870 145.720 167.250 146.725 ;
        RECT 168.090 145.720 170.470 146.725 ;
        RECT 171.310 145.720 173.690 146.725 ;
        RECT 174.530 145.720 176.910 146.725 ;
        RECT 177.750 145.720 180.130 146.725 ;
        RECT 180.970 145.720 183.350 146.725 ;
        RECT 184.190 145.720 186.570 146.725 ;
        RECT 187.410 145.720 189.790 146.725 ;
        RECT 190.630 145.720 193.010 146.725 ;
        RECT 193.850 145.720 196.230 146.725 ;
        RECT 197.070 145.720 202.670 146.725 ;
        RECT 203.510 145.720 205.890 146.725 ;
        RECT 206.730 145.720 209.110 146.725 ;
        RECT 209.950 145.720 212.330 146.725 ;
        RECT 213.170 145.720 215.550 146.725 ;
        RECT 216.390 145.720 218.770 146.725 ;
        RECT 219.610 145.720 221.990 146.725 ;
        RECT 222.830 145.720 225.210 146.725 ;
        RECT 226.050 145.720 228.430 146.725 ;
        RECT 229.270 145.720 231.650 146.725 ;
        RECT 232.490 145.720 234.870 146.725 ;
        RECT 235.710 145.720 241.310 146.725 ;
        RECT 242.150 145.720 244.530 146.725 ;
        RECT 245.370 145.720 247.750 146.725 ;
        RECT 248.590 145.720 250.970 146.725 ;
        RECT 251.810 145.720 254.190 146.725 ;
        RECT 255.030 145.720 257.410 146.725 ;
        RECT 258.250 145.720 260.630 146.725 ;
        RECT 261.470 145.720 263.850 146.725 ;
        RECT 264.690 145.720 267.070 146.725 ;
        RECT 267.910 145.720 270.290 146.725 ;
        RECT 271.130 145.720 273.510 146.725 ;
        RECT 274.350 145.720 279.950 146.725 ;
        RECT 280.790 145.720 283.170 146.725 ;
        RECT 284.010 145.720 286.390 146.725 ;
        RECT 287.230 145.720 289.610 146.725 ;
        RECT 290.450 145.720 292.830 146.725 ;
        RECT 293.670 145.720 296.050 146.725 ;
        RECT 296.890 145.720 299.270 146.725 ;
        RECT 300.110 145.720 302.490 146.725 ;
        RECT 303.330 145.720 305.710 146.725 ;
        RECT 306.550 145.720 308.930 146.725 ;
        RECT 309.770 145.720 312.150 146.725 ;
        RECT 312.990 145.720 318.590 146.725 ;
        RECT 319.430 145.720 321.810 146.725 ;
        RECT 322.650 145.720 325.030 146.725 ;
        RECT 325.870 145.720 328.250 146.725 ;
        RECT 329.090 145.720 331.470 146.725 ;
        RECT 332.310 145.720 334.690 146.725 ;
        RECT 335.530 145.720 337.910 146.725 ;
        RECT 338.750 145.720 341.130 146.725 ;
        RECT 341.970 145.720 344.350 146.725 ;
        RECT 345.190 145.720 347.570 146.725 ;
        RECT 348.410 145.720 350.790 146.725 ;
        RECT 351.630 145.720 357.230 146.725 ;
        RECT 358.070 145.720 360.450 146.725 ;
        RECT 361.290 145.720 363.670 146.725 ;
        RECT 364.510 145.720 366.890 146.725 ;
        RECT 367.730 145.720 370.110 146.725 ;
        RECT 370.950 145.720 373.330 146.725 ;
        RECT 374.170 145.720 376.550 146.725 ;
        RECT 377.390 145.720 379.770 146.725 ;
        RECT 380.610 145.720 382.990 146.725 ;
        RECT 383.830 145.720 386.210 146.725 ;
        RECT 387.050 145.720 389.430 146.725 ;
        RECT 390.270 145.720 395.870 146.725 ;
        RECT 396.710 145.720 399.090 146.725 ;
        RECT 399.930 145.720 402.310 146.725 ;
        RECT 403.150 145.720 405.530 146.725 ;
        RECT 406.370 145.720 408.750 146.725 ;
        RECT 409.590 145.720 411.970 146.725 ;
        RECT 412.810 145.720 415.190 146.725 ;
        RECT 416.030 145.720 418.410 146.725 ;
        RECT 419.250 145.720 421.630 146.725 ;
        RECT 422.470 145.720 424.850 146.725 ;
        RECT 425.690 145.720 428.070 146.725 ;
        RECT 428.910 145.720 434.510 146.725 ;
        RECT 435.350 145.720 437.730 146.725 ;
        RECT 438.570 145.720 440.950 146.725 ;
        RECT 441.790 145.720 444.170 146.725 ;
        RECT 445.010 145.720 447.390 146.725 ;
        RECT 0.100 4.280 447.940 145.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
        RECT 119.790 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 141.490 4.280 ;
        RECT 142.330 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.930 4.280 ;
        RECT 148.770 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 160.810 4.280 ;
        RECT 161.650 0.155 164.030 4.280 ;
        RECT 164.870 0.155 167.250 4.280 ;
        RECT 168.090 0.155 170.470 4.280 ;
        RECT 171.310 0.155 173.690 4.280 ;
        RECT 174.530 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 186.570 4.280 ;
        RECT 187.410 0.155 193.010 4.280 ;
        RECT 193.850 0.155 196.230 4.280 ;
        RECT 197.070 0.155 199.450 4.280 ;
        RECT 200.290 0.155 202.670 4.280 ;
        RECT 203.510 0.155 205.890 4.280 ;
        RECT 206.730 0.155 209.110 4.280 ;
        RECT 209.950 0.155 212.330 4.280 ;
        RECT 213.170 0.155 215.550 4.280 ;
        RECT 216.390 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.990 4.280 ;
        RECT 222.830 0.155 225.210 4.280 ;
        RECT 226.050 0.155 231.650 4.280 ;
        RECT 232.490 0.155 234.870 4.280 ;
        RECT 235.710 0.155 238.090 4.280 ;
        RECT 238.930 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 247.750 4.280 ;
        RECT 248.590 0.155 250.970 4.280 ;
        RECT 251.810 0.155 254.190 4.280 ;
        RECT 255.030 0.155 257.410 4.280 ;
        RECT 258.250 0.155 260.630 4.280 ;
        RECT 261.470 0.155 263.850 4.280 ;
        RECT 264.690 0.155 270.290 4.280 ;
        RECT 271.130 0.155 273.510 4.280 ;
        RECT 274.350 0.155 276.730 4.280 ;
        RECT 277.570 0.155 279.950 4.280 ;
        RECT 280.790 0.155 283.170 4.280 ;
        RECT 284.010 0.155 286.390 4.280 ;
        RECT 287.230 0.155 289.610 4.280 ;
        RECT 290.450 0.155 292.830 4.280 ;
        RECT 293.670 0.155 296.050 4.280 ;
        RECT 296.890 0.155 299.270 4.280 ;
        RECT 300.110 0.155 305.710 4.280 ;
        RECT 306.550 0.155 308.930 4.280 ;
        RECT 309.770 0.155 312.150 4.280 ;
        RECT 312.990 0.155 315.370 4.280 ;
        RECT 316.210 0.155 318.590 4.280 ;
        RECT 319.430 0.155 321.810 4.280 ;
        RECT 322.650 0.155 325.030 4.280 ;
        RECT 325.870 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.470 4.280 ;
        RECT 332.310 0.155 334.690 4.280 ;
        RECT 335.530 0.155 337.910 4.280 ;
        RECT 338.750 0.155 344.350 4.280 ;
        RECT 345.190 0.155 347.570 4.280 ;
        RECT 348.410 0.155 350.790 4.280 ;
        RECT 351.630 0.155 354.010 4.280 ;
        RECT 354.850 0.155 357.230 4.280 ;
        RECT 358.070 0.155 360.450 4.280 ;
        RECT 361.290 0.155 363.670 4.280 ;
        RECT 364.510 0.155 366.890 4.280 ;
        RECT 367.730 0.155 370.110 4.280 ;
        RECT 370.950 0.155 373.330 4.280 ;
        RECT 374.170 0.155 376.550 4.280 ;
        RECT 377.390 0.155 382.990 4.280 ;
        RECT 383.830 0.155 386.210 4.280 ;
        RECT 387.050 0.155 389.430 4.280 ;
        RECT 390.270 0.155 392.650 4.280 ;
        RECT 393.490 0.155 395.870 4.280 ;
        RECT 396.710 0.155 399.090 4.280 ;
        RECT 399.930 0.155 402.310 4.280 ;
        RECT 403.150 0.155 405.530 4.280 ;
        RECT 406.370 0.155 408.750 4.280 ;
        RECT 409.590 0.155 411.970 4.280 ;
        RECT 412.810 0.155 415.190 4.280 ;
        RECT 416.030 0.155 421.630 4.280 ;
        RECT 422.470 0.155 424.850 4.280 ;
        RECT 425.690 0.155 428.070 4.280 ;
        RECT 428.910 0.155 431.290 4.280 ;
        RECT 432.130 0.155 434.510 4.280 ;
        RECT 435.350 0.155 437.730 4.280 ;
        RECT 438.570 0.155 440.950 4.280 ;
        RECT 441.790 0.155 444.170 4.280 ;
        RECT 445.010 0.155 447.390 4.280 ;
      LAYER met3 ;
        RECT 4.400 145.840 445.600 146.705 ;
        RECT 4.000 143.840 446.000 145.840 ;
        RECT 4.400 142.440 445.600 143.840 ;
        RECT 4.000 140.440 446.000 142.440 ;
        RECT 4.400 139.040 445.600 140.440 ;
        RECT 4.000 137.040 446.000 139.040 ;
        RECT 4.400 135.640 445.600 137.040 ;
        RECT 4.000 133.640 446.000 135.640 ;
        RECT 4.400 132.240 445.600 133.640 ;
        RECT 4.000 130.240 446.000 132.240 ;
        RECT 4.400 128.840 446.000 130.240 ;
        RECT 4.000 126.840 446.000 128.840 ;
        RECT 4.400 125.440 445.600 126.840 ;
        RECT 4.000 123.440 446.000 125.440 ;
        RECT 4.400 122.040 445.600 123.440 ;
        RECT 4.000 120.040 446.000 122.040 ;
        RECT 4.000 118.640 445.600 120.040 ;
        RECT 4.000 116.640 446.000 118.640 ;
        RECT 4.400 115.240 445.600 116.640 ;
        RECT 4.000 113.240 446.000 115.240 ;
        RECT 4.400 111.840 445.600 113.240 ;
        RECT 4.000 109.840 446.000 111.840 ;
        RECT 4.400 108.440 445.600 109.840 ;
        RECT 4.000 106.440 446.000 108.440 ;
        RECT 4.400 105.040 445.600 106.440 ;
        RECT 4.000 103.040 446.000 105.040 ;
        RECT 4.400 101.640 445.600 103.040 ;
        RECT 4.000 99.640 446.000 101.640 ;
        RECT 4.400 98.240 445.600 99.640 ;
        RECT 4.000 96.240 446.000 98.240 ;
        RECT 4.400 94.840 445.600 96.240 ;
        RECT 4.000 92.840 446.000 94.840 ;
        RECT 4.400 91.440 445.600 92.840 ;
        RECT 4.000 89.440 446.000 91.440 ;
        RECT 4.400 88.040 446.000 89.440 ;
        RECT 4.000 86.040 446.000 88.040 ;
        RECT 4.400 84.640 445.600 86.040 ;
        RECT 4.000 82.640 446.000 84.640 ;
        RECT 4.400 81.240 445.600 82.640 ;
        RECT 4.000 79.240 446.000 81.240 ;
        RECT 4.000 77.840 445.600 79.240 ;
        RECT 4.000 75.840 446.000 77.840 ;
        RECT 4.400 74.440 445.600 75.840 ;
        RECT 4.000 72.440 446.000 74.440 ;
        RECT 4.400 71.040 445.600 72.440 ;
        RECT 4.000 69.040 446.000 71.040 ;
        RECT 4.400 67.640 445.600 69.040 ;
        RECT 4.000 65.640 446.000 67.640 ;
        RECT 4.400 64.240 445.600 65.640 ;
        RECT 4.000 62.240 446.000 64.240 ;
        RECT 4.400 60.840 445.600 62.240 ;
        RECT 4.000 58.840 446.000 60.840 ;
        RECT 4.400 57.440 445.600 58.840 ;
        RECT 4.000 55.440 446.000 57.440 ;
        RECT 4.400 54.040 445.600 55.440 ;
        RECT 4.000 52.040 446.000 54.040 ;
        RECT 4.400 50.640 445.600 52.040 ;
        RECT 4.000 48.640 446.000 50.640 ;
        RECT 4.400 47.240 446.000 48.640 ;
        RECT 4.000 45.240 446.000 47.240 ;
        RECT 4.400 43.840 445.600 45.240 ;
        RECT 4.000 41.840 446.000 43.840 ;
        RECT 4.400 40.440 445.600 41.840 ;
        RECT 4.000 38.440 446.000 40.440 ;
        RECT 4.000 37.040 445.600 38.440 ;
        RECT 4.000 35.040 446.000 37.040 ;
        RECT 4.400 33.640 445.600 35.040 ;
        RECT 4.000 31.640 446.000 33.640 ;
        RECT 4.400 30.240 445.600 31.640 ;
        RECT 4.000 28.240 446.000 30.240 ;
        RECT 4.400 26.840 445.600 28.240 ;
        RECT 4.000 24.840 446.000 26.840 ;
        RECT 4.400 23.440 445.600 24.840 ;
        RECT 4.000 21.440 446.000 23.440 ;
        RECT 4.400 20.040 445.600 21.440 ;
        RECT 4.000 18.040 446.000 20.040 ;
        RECT 4.400 16.640 445.600 18.040 ;
        RECT 4.000 14.640 446.000 16.640 ;
        RECT 4.400 13.240 445.600 14.640 ;
        RECT 4.000 11.240 446.000 13.240 ;
        RECT 4.400 9.840 445.600 11.240 ;
        RECT 4.000 7.840 446.000 9.840 ;
        RECT 4.400 6.440 446.000 7.840 ;
        RECT 4.000 4.440 446.000 6.440 ;
        RECT 4.400 3.040 445.600 4.440 ;
        RECT 4.000 1.040 446.000 3.040 ;
        RECT 4.000 0.175 445.600 1.040 ;
      LAYER met4 ;
        RECT 132.775 51.175 168.930 129.025 ;
        RECT 171.330 51.175 223.800 129.025 ;
        RECT 226.200 51.175 278.670 129.025 ;
        RECT 281.070 51.175 321.705 129.025 ;
  END
END l1icache_32
END LIBRARY

