VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core_empty
  CLASS BLOCK ;
  FOREIGN core_empty ;
  ORIGIN 0.000 0.000 ;
  SIZE 1600.000 BY 1600.000 ;
  PIN back2dcache_lsq_index_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END back2dcache_lsq_index_o
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 1596.000 1275.490 1600.000 ;
    END
  END clk
  PIN dcache2back_resp_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 1596.000 451.170 1600.000 ;
    END
  END dcache2back_resp_data_i[0]
  PIN dcache2back_resp_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1275.040 1600.000 1275.640 ;
    END
  END dcache2back_resp_data_i[10]
  PIN dcache2back_resp_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 0.000 1372.090 4.000 ;
    END
  END dcache2back_resp_data_i[11]
  PIN dcache2back_resp_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1346.440 1600.000 1347.040 ;
    END
  END dcache2back_resp_data_i[12]
  PIN dcache2back_resp_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END dcache2back_resp_data_i[13]
  PIN dcache2back_resp_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 1596.000 1062.970 1600.000 ;
    END
  END dcache2back_resp_data_i[14]
  PIN dcache2back_resp_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 1596.000 267.630 1600.000 ;
    END
  END dcache2back_resp_data_i[15]
  PIN dcache2back_resp_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 1596.000 567.090 1600.000 ;
    END
  END dcache2back_resp_data_i[16]
  PIN dcache2back_resp_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END dcache2back_resp_data_i[17]
  PIN dcache2back_resp_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1033.640 1600.000 1034.240 ;
    END
  END dcache2back_resp_data_i[18]
  PIN dcache2back_resp_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END dcache2back_resp_data_i[19]
  PIN dcache2back_resp_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END dcache2back_resp_data_i[1]
  PIN dcache2back_resp_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END dcache2back_resp_data_i[20]
  PIN dcache2back_resp_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END dcache2back_resp_data_i[21]
  PIN dcache2back_resp_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END dcache2back_resp_data_i[22]
  PIN dcache2back_resp_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 1596.000 1523.430 1600.000 ;
    END
  END dcache2back_resp_data_i[23]
  PIN dcache2back_resp_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END dcache2back_resp_data_i[24]
  PIN dcache2back_resp_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 1596.000 947.050 1600.000 ;
    END
  END dcache2back_resp_data_i[25]
  PIN dcache2back_resp_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1203.640 4.000 1204.240 ;
    END
  END dcache2back_resp_data_i[26]
  PIN dcache2back_resp_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 1596.000 415.750 1600.000 ;
    END
  END dcache2back_resp_data_i[27]
  PIN dcache2back_resp_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 105.440 1600.000 106.040 ;
    END
  END dcache2back_resp_data_i[28]
  PIN dcache2back_resp_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END dcache2back_resp_data_i[29]
  PIN dcache2back_resp_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END dcache2back_resp_data_i[2]
  PIN dcache2back_resp_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1570.840 4.000 1571.440 ;
    END
  END dcache2back_resp_data_i[30]
  PIN dcache2back_resp_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 1596.000 1459.030 1600.000 ;
    END
  END dcache2back_resp_data_i[31]
  PIN dcache2back_resp_data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END dcache2back_resp_data_i[32]
  PIN dcache2back_resp_data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 1596.000 1491.230 1600.000 ;
    END
  END dcache2back_resp_data_i[33]
  PIN dcache2back_resp_data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1013.240 1600.000 1013.840 ;
    END
  END dcache2back_resp_data_i[34]
  PIN dcache2back_resp_data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 1596.000 1375.310 1600.000 ;
    END
  END dcache2back_resp_data_i[35]
  PIN dcache2back_resp_data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 1596.000 979.250 1600.000 ;
    END
  END dcache2back_resp_data_i[36]
  PIN dcache2back_resp_data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 1596.000 911.630 1600.000 ;
    END
  END dcache2back_resp_data_i[37]
  PIN dcache2back_resp_data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END dcache2back_resp_data_i[38]
  PIN dcache2back_resp_data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END dcache2back_resp_data_i[39]
  PIN dcache2back_resp_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1540.240 1600.000 1540.840 ;
    END
  END dcache2back_resp_data_i[3]
  PIN dcache2back_resp_data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1156.040 1600.000 1156.640 ;
    END
  END dcache2back_resp_data_i[40]
  PIN dcache2back_resp_data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1596.000 103.410 1600.000 ;
    END
  END dcache2back_resp_data_i[41]
  PIN dcache2back_resp_data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 894.240 1600.000 894.840 ;
    END
  END dcache2back_resp_data_i[42]
  PIN dcache2back_resp_data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END dcache2back_resp_data_i[43]
  PIN dcache2back_resp_data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1596.000 167.810 1600.000 ;
    END
  END dcache2back_resp_data_i[44]
  PIN dcache2back_resp_data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END dcache2back_resp_data_i[45]
  PIN dcache2back_resp_data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1596.000 135.610 1600.000 ;
    END
  END dcache2back_resp_data_i[46]
  PIN dcache2back_resp_data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END dcache2back_resp_data_i[47]
  PIN dcache2back_resp_data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END dcache2back_resp_data_i[48]
  PIN dcache2back_resp_data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 1596.000 219.330 1600.000 ;
    END
  END dcache2back_resp_data_i[49]
  PIN dcache2back_resp_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 0.000 1504.110 4.000 ;
    END
  END dcache2back_resp_data_i[4]
  PIN dcache2back_resp_data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 0.000 1172.450 4.000 ;
    END
  END dcache2back_resp_data_i[50]
  PIN dcache2back_resp_data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 0.000 1320.570 4.000 ;
    END
  END dcache2back_resp_data_i[51]
  PIN dcache2back_resp_data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END dcache2back_resp_data_i[52]
  PIN dcache2back_resp_data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 0.000 1488.010 4.000 ;
    END
  END dcache2back_resp_data_i[53]
  PIN dcache2back_resp_data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 316.240 1600.000 316.840 ;
    END
  END dcache2back_resp_data_i[54]
  PIN dcache2back_resp_data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 0.000 1336.670 4.000 ;
    END
  END dcache2back_resp_data_i[55]
  PIN dcache2back_resp_data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END dcache2back_resp_data_i[56]
  PIN dcache2back_resp_data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 1596.000 1211.090 1600.000 ;
    END
  END dcache2back_resp_data_i[57]
  PIN dcache2back_resp_data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 1596.000 547.770 1600.000 ;
    END
  END dcache2back_resp_data_i[58]
  PIN dcache2back_resp_data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1468.840 1600.000 1469.440 ;
    END
  END dcache2back_resp_data_i[59]
  PIN dcache2back_resp_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1557.240 1600.000 1557.840 ;
    END
  END dcache2back_resp_data_i[5]
  PIN dcache2back_resp_data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 612.040 1600.000 612.640 ;
    END
  END dcache2back_resp_data_i[60]
  PIN dcache2back_resp_data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1258.040 1600.000 1258.640 ;
    END
  END dcache2back_resp_data_i[61]
  PIN dcache2back_resp_data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 1596.000 1159.570 1600.000 ;
    END
  END dcache2back_resp_data_i[62]
  PIN dcache2back_resp_data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1533.440 4.000 1534.040 ;
    END
  END dcache2back_resp_data_i[63]
  PIN dcache2back_resp_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 629.040 1600.000 629.640 ;
    END
  END dcache2back_resp_data_i[6]
  PIN dcache2back_resp_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1380.440 1600.000 1381.040 ;
    END
  END dcache2back_resp_data_i[7]
  PIN dcache2back_resp_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1596.000 251.530 1600.000 ;
    END
  END dcache2back_resp_data_i[8]
  PIN dcache2back_resp_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 1596.000 431.850 1600.000 ;
    END
  END dcache2back_resp_data_i[9]
  PIN dcache2back_resp_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1241.040 1600.000 1241.640 ;
    END
  END dcache2back_resp_valid_i
  PIN dcache2back_rob_index_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1596.000 399.650 1600.000 ;
    END
  END dcache2back_rob_index_i
  PIN dcache_opcode
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END dcache_opcode
  PIN dcache_req_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 1596.000 1095.170 1600.000 ;
    END
  END dcache_req_addr[0]
  PIN dcache_req_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 159.840 1600.000 160.440 ;
    END
  END dcache_req_addr[10]
  PIN dcache_req_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END dcache_req_addr[11]
  PIN dcache_req_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1186.640 4.000 1187.240 ;
    END
  END dcache_req_addr[12]
  PIN dcache_req_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1499.440 4.000 1500.040 ;
    END
  END dcache_req_addr[13]
  PIN dcache_req_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1596.000 747.410 1600.000 ;
    END
  END dcache_req_addr[14]
  PIN dcache_req_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 822.840 1600.000 823.440 ;
    END
  END dcache_req_addr[15]
  PIN dcache_req_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1237.640 4.000 1238.240 ;
    END
  END dcache_req_addr[16]
  PIN dcache_req_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 210.840 1600.000 211.440 ;
    END
  END dcache_req_addr[17]
  PIN dcache_req_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 0.000 1404.290 4.000 ;
    END
  END dcache_req_addr[18]
  PIN dcache_req_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END dcache_req_addr[19]
  PIN dcache_req_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1169.640 4.000 1170.240 ;
    END
  END dcache_req_addr[1]
  PIN dcache_req_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END dcache_req_addr[20]
  PIN dcache_req_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 71.440 1600.000 72.040 ;
    END
  END dcache_req_addr[21]
  PIN dcache_req_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 527.040 1600.000 527.640 ;
    END
  END dcache_req_addr[22]
  PIN dcache_req_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 1596.000 383.550 1600.000 ;
    END
  END dcache_req_addr[23]
  PIN dcache_req_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END dcache_req_addr[24]
  PIN dcache_req_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 1596.000 895.530 1600.000 ;
    END
  END dcache_req_addr[25]
  PIN dcache_req_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 0.000 1436.490 4.000 ;
    END
  END dcache_req_addr[26]
  PIN dcache_req_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 299.240 1600.000 299.840 ;
    END
  END dcache_req_addr[27]
  PIN dcache_req_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 1596.000 467.270 1600.000 ;
    END
  END dcache_req_addr[28]
  PIN dcache_req_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END dcache_req_addr[29]
  PIN dcache_req_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END dcache_req_addr[2]
  PIN dcache_req_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 1596.000 847.230 1600.000 ;
    END
  END dcache_req_addr[30]
  PIN dcache_req_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END dcache_req_addr[31]
  PIN dcache_req_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 0.000 1568.510 4.000 ;
    END
  END dcache_req_addr[3]
  PIN dcache_req_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1084.640 1600.000 1085.240 ;
    END
  END dcache_req_addr[4]
  PIN dcache_req_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 1596.000 1442.930 1600.000 ;
    END
  END dcache_req_addr[5]
  PIN dcache_req_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 996.240 1600.000 996.840 ;
    END
  END dcache_req_addr[6]
  PIN dcache_req_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1295.440 1600.000 1296.040 ;
    END
  END dcache_req_addr[7]
  PIN dcache_req_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END dcache_req_addr[8]
  PIN dcache_req_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 1596.000 151.710 1600.000 ;
    END
  END dcache_req_addr[9]
  PIN dcache_req_ready_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END dcache_req_ready_i
  PIN dcache_req_valid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 1596.000 699.110 1600.000 ;
    END
  END dcache_req_valid_o
  PIN dcache_resp_ready_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1596.000 67.990 1600.000 ;
    END
  END dcache_resp_ready_o
  PIN dcache_st_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 510.040 1600.000 510.640 ;
    END
  END dcache_st_data_o[0]
  PIN dcache_st_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END dcache_st_data_o[10]
  PIN dcache_st_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END dcache_st_data_o[11]
  PIN dcache_st_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END dcache_st_data_o[12]
  PIN dcache_st_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 472.640 1600.000 473.240 ;
    END
  END dcache_st_data_o[13]
  PIN dcache_st_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 962.240 1600.000 962.840 ;
    END
  END dcache_st_data_o[14]
  PIN dcache_st_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END dcache_st_data_o[15]
  PIN dcache_st_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END dcache_st_data_o[16]
  PIN dcache_st_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END dcache_st_data_o[17]
  PIN dcache_st_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1485.840 1600.000 1486.440 ;
    END
  END dcache_st_data_o[18]
  PIN dcache_st_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 1596.000 1111.270 1600.000 ;
    END
  END dcache_st_data_o[19]
  PIN dcache_st_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 4.000 ;
    END
  END dcache_st_data_o[1]
  PIN dcache_st_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 1596.000 3.590 1600.000 ;
    END
  END dcache_st_data_o[20]
  PIN dcache_st_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END dcache_st_data_o[21]
  PIN dcache_st_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END dcache_st_data_o[22]
  PIN dcache_st_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 1596.000 1407.510 1600.000 ;
    END
  END dcache_st_data_o[23]
  PIN dcache_st_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 751.440 1600.000 752.040 ;
    END
  END dcache_st_data_o[24]
  PIN dcache_st_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END dcache_st_data_o[25]
  PIN dcache_st_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 142.840 1600.000 143.440 ;
    END
  END dcache_st_data_o[26]
  PIN dcache_st_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END dcache_st_data_o[27]
  PIN dcache_st_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 88.440 1600.000 89.040 ;
    END
  END dcache_st_data_o[28]
  PIN dcache_st_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END dcache_st_data_o[29]
  PIN dcache_st_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1312.440 1600.000 1313.040 ;
    END
  END dcache_st_data_o[2]
  PIN dcache_st_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 1596.000 1011.450 1600.000 ;
    END
  END dcache_st_data_o[30]
  PIN dcache_st_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.040 4.000 1309.640 ;
    END
  END dcache_st_data_o[31]
  PIN dcache_st_data_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END dcache_st_data_o[32]
  PIN dcache_st_data_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END dcache_st_data_o[33]
  PIN dcache_st_data_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 387.640 1600.000 388.240 ;
    END
  END dcache_st_data_o[34]
  PIN dcache_st_data_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END dcache_st_data_o[35]
  PIN dcache_st_data_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END dcache_st_data_o[36]
  PIN dcache_st_data_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END dcache_st_data_o[37]
  PIN dcache_st_data_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END dcache_st_data_o[38]
  PIN dcache_st_data_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 227.840 1600.000 228.440 ;
    END
  END dcache_st_data_o[39]
  PIN dcache_st_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 1596.000 1343.110 1600.000 ;
    END
  END dcache_st_data_o[3]
  PIN dcache_st_data_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.840 4.000 1554.440 ;
    END
  END dcache_st_data_o[40]
  PIN dcache_st_data_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 1596.000 963.150 1600.000 ;
    END
  END dcache_st_data_o[41]
  PIN dcache_st_data_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 489.640 1600.000 490.240 ;
    END
  END dcache_st_data_o[42]
  PIN dcache_st_data_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END dcache_st_data_o[43]
  PIN dcache_st_data_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END dcache_st_data_o[44]
  PIN dcache_st_data_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END dcache_st_data_o[45]
  PIN dcache_st_data_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 333.240 1600.000 333.840 ;
    END
  END dcache_st_data_o[46]
  PIN dcache_st_data_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END dcache_st_data_o[47]
  PIN dcache_st_data_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 544.040 1600.000 544.640 ;
    END
  END dcache_st_data_o[48]
  PIN dcache_st_data_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END dcache_st_data_o[49]
  PIN dcache_st_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 945.240 1600.000 945.840 ;
    END
  END dcache_st_data_o[4]
  PIN dcache_st_data_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.770 1596.000 1591.050 1600.000 ;
    END
  END dcache_st_data_o[50]
  PIN dcache_st_data_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 438.640 1600.000 439.240 ;
    END
  END dcache_st_data_o[51]
  PIN dcache_st_data_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1363.440 1600.000 1364.040 ;
    END
  END dcache_st_data_o[52]
  PIN dcache_st_data_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 788.840 1600.000 789.440 ;
    END
  END dcache_st_data_o[53]
  PIN dcache_st_data_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 1596.000 1027.550 1600.000 ;
    END
  END dcache_st_data_o[54]
  PIN dcache_st_data_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END dcache_st_data_o[55]
  PIN dcache_st_data_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 193.840 1600.000 194.440 ;
    END
  END dcache_st_data_o[56]
  PIN dcache_st_data_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 1596.000 930.950 1600.000 ;
    END
  END dcache_st_data_o[57]
  PIN dcache_st_data_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END dcache_st_data_o[58]
  PIN dcache_st_data_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END dcache_st_data_o[59]
  PIN dcache_st_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 1596.000 631.490 1600.000 ;
    END
  END dcache_st_data_o[5]
  PIN dcache_st_data_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END dcache_st_data_o[60]
  PIN dcache_st_data_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END dcache_st_data_o[61]
  PIN dcache_st_data_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END dcache_st_data_o[62]
  PIN dcache_st_data_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1596.000 19.690 1600.000 ;
    END
  END dcache_st_data_o[63]
  PIN dcache_st_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END dcache_st_data_o[6]
  PIN dcache_st_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 1596.000 795.710 1600.000 ;
    END
  END dcache_st_data_o[7]
  PIN dcache_st_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END dcache_st_data_o[8]
  PIN dcache_st_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 1596.000 1475.130 1600.000 ;
    END
  END dcache_st_data_o[9]
  PIN dcache_type_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1596.000 87.310 1600.000 ;
    END
  END dcache_type_o[0]
  PIN dcache_type_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 367.240 1600.000 367.840 ;
    END
  END dcache_type_o[1]
  PIN dcache_type_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 1596.000 335.250 1600.000 ;
    END
  END dcache_type_o[2]
  PIN icache_req_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1519.840 1600.000 1520.440 ;
    END
  END icache_req_addr[0]
  PIN icache_req_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END icache_req_addr[10]
  PIN icache_req_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END icache_req_addr[11]
  PIN icache_req_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 248.240 1600.000 248.840 ;
    END
  END icache_req_addr[12]
  PIN icache_req_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1050.640 1600.000 1051.240 ;
    END
  END icache_req_addr[13]
  PIN icache_req_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END icache_req_addr[14]
  PIN icache_req_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END icache_req_addr[15]
  PIN icache_req_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END icache_req_addr[16]
  PIN icache_req_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END icache_req_addr[17]
  PIN icache_req_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1292.040 4.000 1292.640 ;
    END
  END icache_req_addr[18]
  PIN icache_req_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 1596.000 1227.190 1600.000 ;
    END
  END icache_req_addr[19]
  PIN icache_req_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END icache_req_addr[1]
  PIN icache_req_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 578.040 1600.000 578.640 ;
    END
  END icache_req_addr[20]
  PIN icache_req_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 1596.000 183.910 1600.000 ;
    END
  END icache_req_addr[21]
  PIN icache_req_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END icache_req_addr[22]
  PIN icache_req_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1271.640 4.000 1272.240 ;
    END
  END icache_req_addr[23]
  PIN icache_req_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END icache_req_addr[24]
  PIN icache_req_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 839.840 1600.000 840.440 ;
    END
  END icache_req_addr[25]
  PIN icache_req_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END icache_req_addr[26]
  PIN icache_req_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1596.000 235.430 1600.000 ;
    END
  END icache_req_addr[27]
  PIN icache_req_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 717.440 1600.000 718.040 ;
    END
  END icache_req_addr[28]
  PIN icache_req_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 4.000 1449.040 ;
    END
  END icache_req_addr[29]
  PIN icache_req_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END icache_req_addr[2]
  PIN icache_req_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 1596.000 1291.590 1600.000 ;
    END
  END icache_req_addr[30]
  PIN icache_req_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1587.840 4.000 1588.440 ;
    END
  END icache_req_addr[31]
  PIN icache_req_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END icache_req_addr[3]
  PIN icache_req_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END icache_req_addr[4]
  PIN icache_req_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1596.000 779.610 1600.000 ;
    END
  END icache_req_addr[5]
  PIN icache_req_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 265.240 1600.000 265.840 ;
    END
  END icache_req_addr[6]
  PIN icache_req_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 1596.000 995.350 1600.000 ;
    END
  END icache_req_addr[7]
  PIN icache_req_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END icache_req_addr[8]
  PIN icache_req_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 561.040 1600.000 561.640 ;
    END
  END icache_req_addr[9]
  PIN icache_req_ready_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1596.000 35.790 1600.000 ;
    END
  END icache_req_ready_i
  PIN icache_req_valid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END icache_req_valid_o
  PIN icache_resp_address_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 1596.000 531.670 1600.000 ;
    END
  END icache_resp_address_i[0]
  PIN icache_resp_address_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 1596.000 663.690 1600.000 ;
    END
  END icache_resp_address_i[10]
  PIN icache_resp_address_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 734.440 1600.000 735.040 ;
    END
  END icache_resp_address_i[11]
  PIN icache_resp_address_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END icache_resp_address_i[12]
  PIN icache_resp_address_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END icache_resp_address_i[13]
  PIN icache_resp_address_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END icache_resp_address_i[14]
  PIN icache_resp_address_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END icache_resp_address_i[15]
  PIN icache_resp_address_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END icache_resp_address_i[16]
  PIN icache_resp_address_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 0.000 1584.610 4.000 ;
    END
  END icache_resp_address_i[17]
  PIN icache_resp_address_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 1596.000 319.150 1600.000 ;
    END
  END icache_resp_address_i[18]
  PIN icache_resp_address_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 1596.000 815.030 1600.000 ;
    END
  END icache_resp_address_i[19]
  PIN icache_resp_address_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1574.240 1600.000 1574.840 ;
    END
  END icache_resp_address_i[1]
  PIN icache_resp_address_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 1596.000 1426.830 1600.000 ;
    END
  END icache_resp_address_i[20]
  PIN icache_resp_address_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END icache_resp_address_i[21]
  PIN icache_resp_address_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 805.840 1600.000 806.440 ;
    END
  END icache_resp_address_i[22]
  PIN icache_resp_address_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 0.000 1304.470 4.000 ;
    END
  END icache_resp_address_i[23]
  PIN icache_resp_address_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END icache_resp_address_i[24]
  PIN icache_resp_address_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END icache_resp_address_i[25]
  PIN icache_resp_address_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 666.440 1600.000 667.040 ;
    END
  END icache_resp_address_i[26]
  PIN icache_resp_address_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1220.640 4.000 1221.240 ;
    END
  END icache_resp_address_i[27]
  PIN icache_resp_address_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1417.840 1600.000 1418.440 ;
    END
  END icache_resp_address_i[28]
  PIN icache_resp_address_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1190.040 1600.000 1190.640 ;
    END
  END icache_resp_address_i[29]
  PIN icache_resp_address_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1135.640 1600.000 1136.240 ;
    END
  END icache_resp_address_i[2]
  PIN icache_resp_address_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1118.640 1600.000 1119.240 ;
    END
  END icache_resp_address_i[30]
  PIN icache_resp_address_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END icache_resp_address_i[31]
  PIN icache_resp_address_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1591.240 1600.000 1591.840 ;
    END
  END icache_resp_address_i[3]
  PIN icache_resp_address_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1596.000 763.510 1600.000 ;
    END
  END icache_resp_address_i[4]
  PIN icache_resp_address_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END icache_resp_address_i[5]
  PIN icache_resp_address_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END icache_resp_address_i[6]
  PIN icache_resp_address_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END icache_resp_address_i[7]
  PIN icache_resp_address_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 0.000 1536.310 4.000 ;
    END
  END icache_resp_address_i[8]
  PIN icache_resp_address_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1502.840 1600.000 1503.440 ;
    END
  END icache_resp_address_i[9]
  PIN icache_resp_ready_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 54.440 1600.000 55.040 ;
    END
  END icache_resp_ready_o
  PIN icache_resp_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 1596.000 831.130 1600.000 ;
    END
  END icache_resp_valid_i
  PIN insn_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END insn_i[0]
  PIN insn_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END insn_i[10]
  PIN insn_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END insn_i[11]
  PIN insn_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1596.000 299.830 1600.000 ;
    END
  END insn_i[12]
  PIN insn_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END insn_i[13]
  PIN insn_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END insn_i[14]
  PIN insn_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END insn_i[15]
  PIN insn_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END insn_i[16]
  PIN insn_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 1596.000 367.450 1600.000 ;
    END
  END insn_i[17]
  PIN insn_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END insn_i[18]
  PIN insn_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 1596.000 731.310 1600.000 ;
    END
  END insn_i[19]
  PIN insn_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 4.000 ;
    END
  END insn_i[1]
  PIN insn_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 1596.000 51.890 1600.000 ;
    END
  END insn_i[20]
  PIN insn_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 1596.000 1259.390 1600.000 ;
    END
  END insn_i[21]
  PIN insn_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 700.440 1600.000 701.040 ;
    END
  END insn_i[22]
  PIN insn_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.040 4.000 1326.640 ;
    END
  END insn_i[23]
  PIN insn_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 1596.000 1558.850 1600.000 ;
    END
  END insn_i[24]
  PIN insn_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 37.440 1600.000 38.040 ;
    END
  END insn_i[25]
  PIN insn_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END insn_i[26]
  PIN insn_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END insn_i[27]
  PIN insn_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 1596.000 599.290 1600.000 ;
    END
  END insn_i[28]
  PIN insn_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END insn_i[29]
  PIN insn_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 683.440 1600.000 684.040 ;
    END
  END insn_i[2]
  PIN insn_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1596.000 119.510 1600.000 ;
    END
  END insn_i[30]
  PIN insn_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END insn_i[31]
  PIN insn_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END insn_i[3]
  PIN insn_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 0.000 1420.390 4.000 ;
    END
  END insn_i[4]
  PIN insn_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 1596.000 647.590 1600.000 ;
    END
  END insn_i[5]
  PIN insn_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 1596.000 1507.330 1600.000 ;
    END
  END insn_i[6]
  PIN insn_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1101.640 1600.000 1102.240 ;
    END
  END insn_i[7]
  PIN insn_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 1596.000 583.190 1600.000 ;
    END
  END insn_i[8]
  PIN insn_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 1596.000 715.210 1600.000 ;
    END
  END insn_i[9]
  PIN meip
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 176.840 1600.000 177.440 ;
    END
  END meip
  PIN others_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END others_wb_ack_i
  PIN others_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END others_wb_adr_o[0]
  PIN others_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END others_wb_adr_o[10]
  PIN others_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 1596.000 879.430 1600.000 ;
    END
  END others_wb_adr_o[11]
  PIN others_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1596.000 283.730 1600.000 ;
    END
  END others_wb_adr_o[12]
  PIN others_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END others_wb_adr_o[13]
  PIN others_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END others_wb_adr_o[14]
  PIN others_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1067.640 1600.000 1068.240 ;
    END
  END others_wb_adr_o[15]
  PIN others_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 979.240 1600.000 979.840 ;
    END
  END others_wb_adr_o[16]
  PIN others_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END others_wb_adr_o[17]
  PIN others_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END others_wb_adr_o[18]
  PIN others_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END others_wb_adr_o[19]
  PIN others_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 0.000 1452.590 4.000 ;
    END
  END others_wb_adr_o[1]
  PIN others_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 1596.000 1143.470 1600.000 ;
    END
  END others_wb_adr_o[20]
  PIN others_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END others_wb_adr_o[21]
  PIN others_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END others_wb_adr_o[22]
  PIN others_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END others_wb_adr_o[23]
  PIN others_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 282.240 1600.000 282.840 ;
    END
  END others_wb_adr_o[24]
  PIN others_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 1596.000 351.350 1600.000 ;
    END
  END others_wb_adr_o[25]
  PIN others_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END others_wb_adr_o[26]
  PIN others_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END others_wb_adr_o[27]
  PIN others_wb_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 1596.000 679.790 1600.000 ;
    END
  END others_wb_adr_o[28]
  PIN others_wb_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 856.840 1600.000 857.440 ;
    END
  END others_wb_adr_o[29]
  PIN others_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1451.840 1600.000 1452.440 ;
    END
  END others_wb_adr_o[2]
  PIN others_wb_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END others_wb_adr_o[30]
  PIN others_wb_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 1596.000 1359.210 1600.000 ;
    END
  END others_wb_adr_o[31]
  PIN others_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 595.040 1600.000 595.640 ;
    END
  END others_wb_adr_o[3]
  PIN others_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END others_wb_adr_o[4]
  PIN others_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 1596.000 1327.010 1600.000 ;
    END
  END others_wb_adr_o[5]
  PIN others_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END others_wb_adr_o[6]
  PIN others_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END others_wb_adr_o[7]
  PIN others_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END others_wb_adr_o[8]
  PIN others_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 0.000 1520.210 4.000 ;
    END
  END others_wb_adr_o[9]
  PIN others_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 350.240 1600.000 350.840 ;
    END
  END others_wb_cyc_o
  PIN others_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1596.000 615.390 1600.000 ;
    END
  END others_wb_dat_i[0]
  PIN others_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1329.440 1600.000 1330.040 ;
    END
  END others_wb_dat_i[10]
  PIN others_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END others_wb_dat_i[11]
  PIN others_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END others_wb_dat_i[12]
  PIN others_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END others_wb_dat_i[13]
  PIN others_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END others_wb_dat_i[14]
  PIN others_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END others_wb_dat_i[15]
  PIN others_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END others_wb_dat_i[16]
  PIN others_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END others_wb_dat_i[17]
  PIN others_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 1596.000 1178.890 1600.000 ;
    END
  END others_wb_dat_i[18]
  PIN others_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 1596.000 1542.750 1600.000 ;
    END
  END others_wb_dat_i[19]
  PIN others_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END others_wb_dat_i[1]
  PIN others_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END others_wb_dat_i[20]
  PIN others_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 911.240 1600.000 911.840 ;
    END
  END others_wb_dat_i[21]
  PIN others_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.670 1596.000 1574.950 1600.000 ;
    END
  END others_wb_dat_i[22]
  PIN others_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END others_wb_dat_i[23]
  PIN others_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1207.040 1600.000 1207.640 ;
    END
  END others_wb_dat_i[24]
  PIN others_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 455.640 1600.000 456.240 ;
    END
  END others_wb_dat_i[25]
  PIN others_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END others_wb_dat_i[26]
  PIN others_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 1596.000 1391.410 1600.000 ;
    END
  END others_wb_dat_i[27]
  PIN others_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 1596.000 483.370 1600.000 ;
    END
  END others_wb_dat_i[28]
  PIN others_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END others_wb_dat_i[29]
  PIN others_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 928.240 1600.000 928.840 ;
    END
  END others_wb_dat_i[2]
  PIN others_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END others_wb_dat_i[30]
  PIN others_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 421.640 1600.000 422.240 ;
    END
  END others_wb_dat_i[31]
  PIN others_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END others_wb_dat_i[3]
  PIN others_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 3.440 1600.000 4.040 ;
    END
  END others_wb_dat_i[4]
  PIN others_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END others_wb_dat_i[5]
  PIN others_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END others_wb_dat_i[6]
  PIN others_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 649.440 1600.000 650.040 ;
    END
  END others_wb_dat_i[7]
  PIN others_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 1596.000 1310.910 1600.000 ;
    END
  END others_wb_dat_i[8]
  PIN others_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1397.440 1600.000 1398.040 ;
    END
  END others_wb_dat_i[9]
  PIN others_wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 20.440 1600.000 21.040 ;
    END
  END others_wb_dat_o[0]
  PIN others_wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END others_wb_dat_o[10]
  PIN others_wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 873.840 1600.000 874.440 ;
    END
  END others_wb_dat_o[11]
  PIN others_wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END others_wb_dat_o[12]
  PIN others_wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1434.840 1600.000 1435.440 ;
    END
  END others_wb_dat_o[13]
  PIN others_wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 1596.000 1243.290 1600.000 ;
    END
  END others_wb_dat_o[14]
  PIN others_wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 125.840 1600.000 126.440 ;
    END
  END others_wb_dat_o[15]
  PIN others_wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 1596.000 1194.990 1600.000 ;
    END
  END others_wb_dat_o[16]
  PIN others_wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END others_wb_dat_o[17]
  PIN others_wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END others_wb_dat_o[18]
  PIN others_wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END others_wb_dat_o[19]
  PIN others_wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END others_wb_dat_o[1]
  PIN others_wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 4.000 ;
    END
  END others_wb_dat_o[20]
  PIN others_wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END others_wb_dat_o[21]
  PIN others_wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END others_wb_dat_o[22]
  PIN others_wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 1596.000 499.470 1600.000 ;
    END
  END others_wb_dat_o[23]
  PIN others_wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END others_wb_dat_o[24]
  PIN others_wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END others_wb_dat_o[25]
  PIN others_wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END others_wb_dat_o[26]
  PIN others_wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 1596.000 863.330 1600.000 ;
    END
  END others_wb_dat_o[27]
  PIN others_wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 1596.000 515.570 1600.000 ;
    END
  END others_wb_dat_o[28]
  PIN others_wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END others_wb_dat_o[29]
  PIN others_wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 1596.000 1127.370 1600.000 ;
    END
  END others_wb_dat_o[2]
  PIN others_wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 404.640 1600.000 405.240 ;
    END
  END others_wb_dat_o[30]
  PIN others_wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END others_wb_dat_o[31]
  PIN others_wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1224.040 1600.000 1224.640 ;
    END
  END others_wb_dat_o[3]
  PIN others_wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END others_wb_dat_o[4]
  PIN others_wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END others_wb_dat_o[5]
  PIN others_wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END others_wb_dat_o[6]
  PIN others_wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1173.040 1600.000 1173.640 ;
    END
  END others_wb_dat_o[7]
  PIN others_wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END others_wb_dat_o[8]
  PIN others_wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 1596.000 1079.070 1600.000 ;
    END
  END others_wb_dat_o[9]
  PIN others_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 1596.000 1043.650 1600.000 ;
    END
  END others_wb_sel_o[0]
  PIN others_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1516.440 4.000 1517.040 ;
    END
  END others_wb_sel_o[1]
  PIN others_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 1596.000 203.230 1600.000 ;
    END
  END others_wb_sel_o[2]
  PIN others_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 4.000 ;
    END
  END others_wb_sel_o[3]
  PIN others_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END others_wb_stb_o
  PIN others_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END others_wb_we_o
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 771.840 1600.000 772.440 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1588.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1588.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1594.360 1588.565 ;
      LAYER met1 ;
        RECT 0.070 6.840 1596.130 1591.840 ;
      LAYER met2 ;
        RECT 0.100 1595.720 3.030 1596.370 ;
        RECT 3.870 1595.720 19.130 1596.370 ;
        RECT 19.970 1595.720 35.230 1596.370 ;
        RECT 36.070 1595.720 51.330 1596.370 ;
        RECT 52.170 1595.720 67.430 1596.370 ;
        RECT 68.270 1595.720 86.750 1596.370 ;
        RECT 87.590 1595.720 102.850 1596.370 ;
        RECT 103.690 1595.720 118.950 1596.370 ;
        RECT 119.790 1595.720 135.050 1596.370 ;
        RECT 135.890 1595.720 151.150 1596.370 ;
        RECT 151.990 1595.720 167.250 1596.370 ;
        RECT 168.090 1595.720 183.350 1596.370 ;
        RECT 184.190 1595.720 202.670 1596.370 ;
        RECT 203.510 1595.720 218.770 1596.370 ;
        RECT 219.610 1595.720 234.870 1596.370 ;
        RECT 235.710 1595.720 250.970 1596.370 ;
        RECT 251.810 1595.720 267.070 1596.370 ;
        RECT 267.910 1595.720 283.170 1596.370 ;
        RECT 284.010 1595.720 299.270 1596.370 ;
        RECT 300.110 1595.720 318.590 1596.370 ;
        RECT 319.430 1595.720 334.690 1596.370 ;
        RECT 335.530 1595.720 350.790 1596.370 ;
        RECT 351.630 1595.720 366.890 1596.370 ;
        RECT 367.730 1595.720 382.990 1596.370 ;
        RECT 383.830 1595.720 399.090 1596.370 ;
        RECT 399.930 1595.720 415.190 1596.370 ;
        RECT 416.030 1595.720 431.290 1596.370 ;
        RECT 432.130 1595.720 450.610 1596.370 ;
        RECT 451.450 1595.720 466.710 1596.370 ;
        RECT 467.550 1595.720 482.810 1596.370 ;
        RECT 483.650 1595.720 498.910 1596.370 ;
        RECT 499.750 1595.720 515.010 1596.370 ;
        RECT 515.850 1595.720 531.110 1596.370 ;
        RECT 531.950 1595.720 547.210 1596.370 ;
        RECT 548.050 1595.720 566.530 1596.370 ;
        RECT 567.370 1595.720 582.630 1596.370 ;
        RECT 583.470 1595.720 598.730 1596.370 ;
        RECT 599.570 1595.720 614.830 1596.370 ;
        RECT 615.670 1595.720 630.930 1596.370 ;
        RECT 631.770 1595.720 647.030 1596.370 ;
        RECT 647.870 1595.720 663.130 1596.370 ;
        RECT 663.970 1595.720 679.230 1596.370 ;
        RECT 680.070 1595.720 698.550 1596.370 ;
        RECT 699.390 1595.720 714.650 1596.370 ;
        RECT 715.490 1595.720 730.750 1596.370 ;
        RECT 731.590 1595.720 746.850 1596.370 ;
        RECT 747.690 1595.720 762.950 1596.370 ;
        RECT 763.790 1595.720 779.050 1596.370 ;
        RECT 779.890 1595.720 795.150 1596.370 ;
        RECT 795.990 1595.720 814.470 1596.370 ;
        RECT 815.310 1595.720 830.570 1596.370 ;
        RECT 831.410 1595.720 846.670 1596.370 ;
        RECT 847.510 1595.720 862.770 1596.370 ;
        RECT 863.610 1595.720 878.870 1596.370 ;
        RECT 879.710 1595.720 894.970 1596.370 ;
        RECT 895.810 1595.720 911.070 1596.370 ;
        RECT 911.910 1595.720 930.390 1596.370 ;
        RECT 931.230 1595.720 946.490 1596.370 ;
        RECT 947.330 1595.720 962.590 1596.370 ;
        RECT 963.430 1595.720 978.690 1596.370 ;
        RECT 979.530 1595.720 994.790 1596.370 ;
        RECT 995.630 1595.720 1010.890 1596.370 ;
        RECT 1011.730 1595.720 1026.990 1596.370 ;
        RECT 1027.830 1595.720 1043.090 1596.370 ;
        RECT 1043.930 1595.720 1062.410 1596.370 ;
        RECT 1063.250 1595.720 1078.510 1596.370 ;
        RECT 1079.350 1595.720 1094.610 1596.370 ;
        RECT 1095.450 1595.720 1110.710 1596.370 ;
        RECT 1111.550 1595.720 1126.810 1596.370 ;
        RECT 1127.650 1595.720 1142.910 1596.370 ;
        RECT 1143.750 1595.720 1159.010 1596.370 ;
        RECT 1159.850 1595.720 1178.330 1596.370 ;
        RECT 1179.170 1595.720 1194.430 1596.370 ;
        RECT 1195.270 1595.720 1210.530 1596.370 ;
        RECT 1211.370 1595.720 1226.630 1596.370 ;
        RECT 1227.470 1595.720 1242.730 1596.370 ;
        RECT 1243.570 1595.720 1258.830 1596.370 ;
        RECT 1259.670 1595.720 1274.930 1596.370 ;
        RECT 1275.770 1595.720 1291.030 1596.370 ;
        RECT 1291.870 1595.720 1310.350 1596.370 ;
        RECT 1311.190 1595.720 1326.450 1596.370 ;
        RECT 1327.290 1595.720 1342.550 1596.370 ;
        RECT 1343.390 1595.720 1358.650 1596.370 ;
        RECT 1359.490 1595.720 1374.750 1596.370 ;
        RECT 1375.590 1595.720 1390.850 1596.370 ;
        RECT 1391.690 1595.720 1406.950 1596.370 ;
        RECT 1407.790 1595.720 1426.270 1596.370 ;
        RECT 1427.110 1595.720 1442.370 1596.370 ;
        RECT 1443.210 1595.720 1458.470 1596.370 ;
        RECT 1459.310 1595.720 1474.570 1596.370 ;
        RECT 1475.410 1595.720 1490.670 1596.370 ;
        RECT 1491.510 1595.720 1506.770 1596.370 ;
        RECT 1507.610 1595.720 1522.870 1596.370 ;
        RECT 1523.710 1595.720 1542.190 1596.370 ;
        RECT 1543.030 1595.720 1558.290 1596.370 ;
        RECT 1559.130 1595.720 1574.390 1596.370 ;
        RECT 1575.230 1595.720 1590.490 1596.370 ;
        RECT 1591.330 1595.720 1596.100 1596.370 ;
        RECT 0.100 4.280 1596.100 1595.720 ;
        RECT 0.650 3.555 15.910 4.280 ;
        RECT 16.750 3.555 32.010 4.280 ;
        RECT 32.850 3.555 48.110 4.280 ;
        RECT 48.950 3.555 64.210 4.280 ;
        RECT 65.050 3.555 80.310 4.280 ;
        RECT 81.150 3.555 96.410 4.280 ;
        RECT 97.250 3.555 112.510 4.280 ;
        RECT 113.350 3.555 131.830 4.280 ;
        RECT 132.670 3.555 147.930 4.280 ;
        RECT 148.770 3.555 164.030 4.280 ;
        RECT 164.870 3.555 180.130 4.280 ;
        RECT 180.970 3.555 196.230 4.280 ;
        RECT 197.070 3.555 212.330 4.280 ;
        RECT 213.170 3.555 228.430 4.280 ;
        RECT 229.270 3.555 247.750 4.280 ;
        RECT 248.590 3.555 263.850 4.280 ;
        RECT 264.690 3.555 279.950 4.280 ;
        RECT 280.790 3.555 296.050 4.280 ;
        RECT 296.890 3.555 312.150 4.280 ;
        RECT 312.990 3.555 328.250 4.280 ;
        RECT 329.090 3.555 344.350 4.280 ;
        RECT 345.190 3.555 360.450 4.280 ;
        RECT 361.290 3.555 379.770 4.280 ;
        RECT 380.610 3.555 395.870 4.280 ;
        RECT 396.710 3.555 411.970 4.280 ;
        RECT 412.810 3.555 428.070 4.280 ;
        RECT 428.910 3.555 444.170 4.280 ;
        RECT 445.010 3.555 460.270 4.280 ;
        RECT 461.110 3.555 476.370 4.280 ;
        RECT 477.210 3.555 495.690 4.280 ;
        RECT 496.530 3.555 511.790 4.280 ;
        RECT 512.630 3.555 527.890 4.280 ;
        RECT 528.730 3.555 543.990 4.280 ;
        RECT 544.830 3.555 560.090 4.280 ;
        RECT 560.930 3.555 576.190 4.280 ;
        RECT 577.030 3.555 592.290 4.280 ;
        RECT 593.130 3.555 611.610 4.280 ;
        RECT 612.450 3.555 627.710 4.280 ;
        RECT 628.550 3.555 643.810 4.280 ;
        RECT 644.650 3.555 659.910 4.280 ;
        RECT 660.750 3.555 676.010 4.280 ;
        RECT 676.850 3.555 692.110 4.280 ;
        RECT 692.950 3.555 708.210 4.280 ;
        RECT 709.050 3.555 724.310 4.280 ;
        RECT 725.150 3.555 743.630 4.280 ;
        RECT 744.470 3.555 759.730 4.280 ;
        RECT 760.570 3.555 775.830 4.280 ;
        RECT 776.670 3.555 791.930 4.280 ;
        RECT 792.770 3.555 808.030 4.280 ;
        RECT 808.870 3.555 824.130 4.280 ;
        RECT 824.970 3.555 840.230 4.280 ;
        RECT 841.070 3.555 859.550 4.280 ;
        RECT 860.390 3.555 875.650 4.280 ;
        RECT 876.490 3.555 891.750 4.280 ;
        RECT 892.590 3.555 907.850 4.280 ;
        RECT 908.690 3.555 923.950 4.280 ;
        RECT 924.790 3.555 940.050 4.280 ;
        RECT 940.890 3.555 956.150 4.280 ;
        RECT 956.990 3.555 972.250 4.280 ;
        RECT 973.090 3.555 991.570 4.280 ;
        RECT 992.410 3.555 1007.670 4.280 ;
        RECT 1008.510 3.555 1023.770 4.280 ;
        RECT 1024.610 3.555 1039.870 4.280 ;
        RECT 1040.710 3.555 1055.970 4.280 ;
        RECT 1056.810 3.555 1072.070 4.280 ;
        RECT 1072.910 3.555 1088.170 4.280 ;
        RECT 1089.010 3.555 1107.490 4.280 ;
        RECT 1108.330 3.555 1123.590 4.280 ;
        RECT 1124.430 3.555 1139.690 4.280 ;
        RECT 1140.530 3.555 1155.790 4.280 ;
        RECT 1156.630 3.555 1171.890 4.280 ;
        RECT 1172.730 3.555 1187.990 4.280 ;
        RECT 1188.830 3.555 1204.090 4.280 ;
        RECT 1204.930 3.555 1223.410 4.280 ;
        RECT 1224.250 3.555 1239.510 4.280 ;
        RECT 1240.350 3.555 1255.610 4.280 ;
        RECT 1256.450 3.555 1271.710 4.280 ;
        RECT 1272.550 3.555 1287.810 4.280 ;
        RECT 1288.650 3.555 1303.910 4.280 ;
        RECT 1304.750 3.555 1320.010 4.280 ;
        RECT 1320.850 3.555 1336.110 4.280 ;
        RECT 1336.950 3.555 1355.430 4.280 ;
        RECT 1356.270 3.555 1371.530 4.280 ;
        RECT 1372.370 3.555 1387.630 4.280 ;
        RECT 1388.470 3.555 1403.730 4.280 ;
        RECT 1404.570 3.555 1419.830 4.280 ;
        RECT 1420.670 3.555 1435.930 4.280 ;
        RECT 1436.770 3.555 1452.030 4.280 ;
        RECT 1452.870 3.555 1471.350 4.280 ;
        RECT 1472.190 3.555 1487.450 4.280 ;
        RECT 1488.290 3.555 1503.550 4.280 ;
        RECT 1504.390 3.555 1519.650 4.280 ;
        RECT 1520.490 3.555 1535.750 4.280 ;
        RECT 1536.590 3.555 1551.850 4.280 ;
        RECT 1552.690 3.555 1567.950 4.280 ;
        RECT 1568.790 3.555 1584.050 4.280 ;
        RECT 1584.890 3.555 1596.100 4.280 ;
      LAYER met3 ;
        RECT 4.000 1590.840 1595.600 1591.705 ;
        RECT 4.000 1588.840 1596.000 1590.840 ;
        RECT 4.400 1587.440 1596.000 1588.840 ;
        RECT 4.000 1575.240 1596.000 1587.440 ;
        RECT 4.000 1573.840 1595.600 1575.240 ;
        RECT 4.000 1571.840 1596.000 1573.840 ;
        RECT 4.400 1570.440 1596.000 1571.840 ;
        RECT 4.000 1558.240 1596.000 1570.440 ;
        RECT 4.000 1556.840 1595.600 1558.240 ;
        RECT 4.000 1554.840 1596.000 1556.840 ;
        RECT 4.400 1553.440 1596.000 1554.840 ;
        RECT 4.000 1541.240 1596.000 1553.440 ;
        RECT 4.000 1539.840 1595.600 1541.240 ;
        RECT 4.000 1534.440 1596.000 1539.840 ;
        RECT 4.400 1533.040 1596.000 1534.440 ;
        RECT 4.000 1520.840 1596.000 1533.040 ;
        RECT 4.000 1519.440 1595.600 1520.840 ;
        RECT 4.000 1517.440 1596.000 1519.440 ;
        RECT 4.400 1516.040 1596.000 1517.440 ;
        RECT 4.000 1503.840 1596.000 1516.040 ;
        RECT 4.000 1502.440 1595.600 1503.840 ;
        RECT 4.000 1500.440 1596.000 1502.440 ;
        RECT 4.400 1499.040 1596.000 1500.440 ;
        RECT 4.000 1486.840 1596.000 1499.040 ;
        RECT 4.000 1485.440 1595.600 1486.840 ;
        RECT 4.000 1483.440 1596.000 1485.440 ;
        RECT 4.400 1482.040 1596.000 1483.440 ;
        RECT 4.000 1469.840 1596.000 1482.040 ;
        RECT 4.000 1468.440 1595.600 1469.840 ;
        RECT 4.000 1466.440 1596.000 1468.440 ;
        RECT 4.400 1465.040 1596.000 1466.440 ;
        RECT 4.000 1452.840 1596.000 1465.040 ;
        RECT 4.000 1451.440 1595.600 1452.840 ;
        RECT 4.000 1449.440 1596.000 1451.440 ;
        RECT 4.400 1448.040 1596.000 1449.440 ;
        RECT 4.000 1435.840 1596.000 1448.040 ;
        RECT 4.000 1434.440 1595.600 1435.840 ;
        RECT 4.000 1432.440 1596.000 1434.440 ;
        RECT 4.400 1431.040 1596.000 1432.440 ;
        RECT 4.000 1418.840 1596.000 1431.040 ;
        RECT 4.000 1417.440 1595.600 1418.840 ;
        RECT 4.000 1412.040 1596.000 1417.440 ;
        RECT 4.400 1410.640 1596.000 1412.040 ;
        RECT 4.000 1398.440 1596.000 1410.640 ;
        RECT 4.000 1397.040 1595.600 1398.440 ;
        RECT 4.000 1395.040 1596.000 1397.040 ;
        RECT 4.400 1393.640 1596.000 1395.040 ;
        RECT 4.000 1381.440 1596.000 1393.640 ;
        RECT 4.000 1380.040 1595.600 1381.440 ;
        RECT 4.000 1378.040 1596.000 1380.040 ;
        RECT 4.400 1376.640 1596.000 1378.040 ;
        RECT 4.000 1364.440 1596.000 1376.640 ;
        RECT 4.000 1363.040 1595.600 1364.440 ;
        RECT 4.000 1361.040 1596.000 1363.040 ;
        RECT 4.400 1359.640 1596.000 1361.040 ;
        RECT 4.000 1347.440 1596.000 1359.640 ;
        RECT 4.000 1346.040 1595.600 1347.440 ;
        RECT 4.000 1344.040 1596.000 1346.040 ;
        RECT 4.400 1342.640 1596.000 1344.040 ;
        RECT 4.000 1330.440 1596.000 1342.640 ;
        RECT 4.000 1329.040 1595.600 1330.440 ;
        RECT 4.000 1327.040 1596.000 1329.040 ;
        RECT 4.400 1325.640 1596.000 1327.040 ;
        RECT 4.000 1313.440 1596.000 1325.640 ;
        RECT 4.000 1312.040 1595.600 1313.440 ;
        RECT 4.000 1310.040 1596.000 1312.040 ;
        RECT 4.400 1308.640 1596.000 1310.040 ;
        RECT 4.000 1296.440 1596.000 1308.640 ;
        RECT 4.000 1295.040 1595.600 1296.440 ;
        RECT 4.000 1293.040 1596.000 1295.040 ;
        RECT 4.400 1291.640 1596.000 1293.040 ;
        RECT 4.000 1276.040 1596.000 1291.640 ;
        RECT 4.000 1274.640 1595.600 1276.040 ;
        RECT 4.000 1272.640 1596.000 1274.640 ;
        RECT 4.400 1271.240 1596.000 1272.640 ;
        RECT 4.000 1259.040 1596.000 1271.240 ;
        RECT 4.000 1257.640 1595.600 1259.040 ;
        RECT 4.000 1255.640 1596.000 1257.640 ;
        RECT 4.400 1254.240 1596.000 1255.640 ;
        RECT 4.000 1242.040 1596.000 1254.240 ;
        RECT 4.000 1240.640 1595.600 1242.040 ;
        RECT 4.000 1238.640 1596.000 1240.640 ;
        RECT 4.400 1237.240 1596.000 1238.640 ;
        RECT 4.000 1225.040 1596.000 1237.240 ;
        RECT 4.000 1223.640 1595.600 1225.040 ;
        RECT 4.000 1221.640 1596.000 1223.640 ;
        RECT 4.400 1220.240 1596.000 1221.640 ;
        RECT 4.000 1208.040 1596.000 1220.240 ;
        RECT 4.000 1206.640 1595.600 1208.040 ;
        RECT 4.000 1204.640 1596.000 1206.640 ;
        RECT 4.400 1203.240 1596.000 1204.640 ;
        RECT 4.000 1191.040 1596.000 1203.240 ;
        RECT 4.000 1189.640 1595.600 1191.040 ;
        RECT 4.000 1187.640 1596.000 1189.640 ;
        RECT 4.400 1186.240 1596.000 1187.640 ;
        RECT 4.000 1174.040 1596.000 1186.240 ;
        RECT 4.000 1172.640 1595.600 1174.040 ;
        RECT 4.000 1170.640 1596.000 1172.640 ;
        RECT 4.400 1169.240 1596.000 1170.640 ;
        RECT 4.000 1157.040 1596.000 1169.240 ;
        RECT 4.000 1155.640 1595.600 1157.040 ;
        RECT 4.000 1150.240 1596.000 1155.640 ;
        RECT 4.400 1148.840 1596.000 1150.240 ;
        RECT 4.000 1136.640 1596.000 1148.840 ;
        RECT 4.000 1135.240 1595.600 1136.640 ;
        RECT 4.000 1133.240 1596.000 1135.240 ;
        RECT 4.400 1131.840 1596.000 1133.240 ;
        RECT 4.000 1119.640 1596.000 1131.840 ;
        RECT 4.000 1118.240 1595.600 1119.640 ;
        RECT 4.000 1116.240 1596.000 1118.240 ;
        RECT 4.400 1114.840 1596.000 1116.240 ;
        RECT 4.000 1102.640 1596.000 1114.840 ;
        RECT 4.000 1101.240 1595.600 1102.640 ;
        RECT 4.000 1099.240 1596.000 1101.240 ;
        RECT 4.400 1097.840 1596.000 1099.240 ;
        RECT 4.000 1085.640 1596.000 1097.840 ;
        RECT 4.000 1084.240 1595.600 1085.640 ;
        RECT 4.000 1082.240 1596.000 1084.240 ;
        RECT 4.400 1080.840 1596.000 1082.240 ;
        RECT 4.000 1068.640 1596.000 1080.840 ;
        RECT 4.000 1067.240 1595.600 1068.640 ;
        RECT 4.000 1065.240 1596.000 1067.240 ;
        RECT 4.400 1063.840 1596.000 1065.240 ;
        RECT 4.000 1051.640 1596.000 1063.840 ;
        RECT 4.000 1050.240 1595.600 1051.640 ;
        RECT 4.000 1048.240 1596.000 1050.240 ;
        RECT 4.400 1046.840 1596.000 1048.240 ;
        RECT 4.000 1034.640 1596.000 1046.840 ;
        RECT 4.000 1033.240 1595.600 1034.640 ;
        RECT 4.000 1027.840 1596.000 1033.240 ;
        RECT 4.400 1026.440 1596.000 1027.840 ;
        RECT 4.000 1014.240 1596.000 1026.440 ;
        RECT 4.000 1012.840 1595.600 1014.240 ;
        RECT 4.000 1010.840 1596.000 1012.840 ;
        RECT 4.400 1009.440 1596.000 1010.840 ;
        RECT 4.000 997.240 1596.000 1009.440 ;
        RECT 4.000 995.840 1595.600 997.240 ;
        RECT 4.000 993.840 1596.000 995.840 ;
        RECT 4.400 992.440 1596.000 993.840 ;
        RECT 4.000 980.240 1596.000 992.440 ;
        RECT 4.000 978.840 1595.600 980.240 ;
        RECT 4.000 976.840 1596.000 978.840 ;
        RECT 4.400 975.440 1596.000 976.840 ;
        RECT 4.000 963.240 1596.000 975.440 ;
        RECT 4.000 961.840 1595.600 963.240 ;
        RECT 4.000 959.840 1596.000 961.840 ;
        RECT 4.400 958.440 1596.000 959.840 ;
        RECT 4.000 946.240 1596.000 958.440 ;
        RECT 4.000 944.840 1595.600 946.240 ;
        RECT 4.000 942.840 1596.000 944.840 ;
        RECT 4.400 941.440 1596.000 942.840 ;
        RECT 4.000 929.240 1596.000 941.440 ;
        RECT 4.000 927.840 1595.600 929.240 ;
        RECT 4.000 925.840 1596.000 927.840 ;
        RECT 4.400 924.440 1596.000 925.840 ;
        RECT 4.000 912.240 1596.000 924.440 ;
        RECT 4.000 910.840 1595.600 912.240 ;
        RECT 4.000 908.840 1596.000 910.840 ;
        RECT 4.400 907.440 1596.000 908.840 ;
        RECT 4.000 895.240 1596.000 907.440 ;
        RECT 4.000 893.840 1595.600 895.240 ;
        RECT 4.000 888.440 1596.000 893.840 ;
        RECT 4.400 887.040 1596.000 888.440 ;
        RECT 4.000 874.840 1596.000 887.040 ;
        RECT 4.000 873.440 1595.600 874.840 ;
        RECT 4.000 871.440 1596.000 873.440 ;
        RECT 4.400 870.040 1596.000 871.440 ;
        RECT 4.000 857.840 1596.000 870.040 ;
        RECT 4.000 856.440 1595.600 857.840 ;
        RECT 4.000 854.440 1596.000 856.440 ;
        RECT 4.400 853.040 1596.000 854.440 ;
        RECT 4.000 840.840 1596.000 853.040 ;
        RECT 4.000 839.440 1595.600 840.840 ;
        RECT 4.000 837.440 1596.000 839.440 ;
        RECT 4.400 836.040 1596.000 837.440 ;
        RECT 4.000 823.840 1596.000 836.040 ;
        RECT 4.000 822.440 1595.600 823.840 ;
        RECT 4.000 820.440 1596.000 822.440 ;
        RECT 4.400 819.040 1596.000 820.440 ;
        RECT 4.000 806.840 1596.000 819.040 ;
        RECT 4.000 805.440 1595.600 806.840 ;
        RECT 4.000 803.440 1596.000 805.440 ;
        RECT 4.400 802.040 1596.000 803.440 ;
        RECT 4.000 789.840 1596.000 802.040 ;
        RECT 4.000 788.440 1595.600 789.840 ;
        RECT 4.000 786.440 1596.000 788.440 ;
        RECT 4.400 785.040 1596.000 786.440 ;
        RECT 4.000 772.840 1596.000 785.040 ;
        RECT 4.000 771.440 1595.600 772.840 ;
        RECT 4.000 766.040 1596.000 771.440 ;
        RECT 4.400 764.640 1596.000 766.040 ;
        RECT 4.000 752.440 1596.000 764.640 ;
        RECT 4.000 751.040 1595.600 752.440 ;
        RECT 4.000 749.040 1596.000 751.040 ;
        RECT 4.400 747.640 1596.000 749.040 ;
        RECT 4.000 735.440 1596.000 747.640 ;
        RECT 4.000 734.040 1595.600 735.440 ;
        RECT 4.000 732.040 1596.000 734.040 ;
        RECT 4.400 730.640 1596.000 732.040 ;
        RECT 4.000 718.440 1596.000 730.640 ;
        RECT 4.000 717.040 1595.600 718.440 ;
        RECT 4.000 715.040 1596.000 717.040 ;
        RECT 4.400 713.640 1596.000 715.040 ;
        RECT 4.000 701.440 1596.000 713.640 ;
        RECT 4.000 700.040 1595.600 701.440 ;
        RECT 4.000 698.040 1596.000 700.040 ;
        RECT 4.400 696.640 1596.000 698.040 ;
        RECT 4.000 684.440 1596.000 696.640 ;
        RECT 4.000 683.040 1595.600 684.440 ;
        RECT 4.000 681.040 1596.000 683.040 ;
        RECT 4.400 679.640 1596.000 681.040 ;
        RECT 4.000 667.440 1596.000 679.640 ;
        RECT 4.000 666.040 1595.600 667.440 ;
        RECT 4.000 664.040 1596.000 666.040 ;
        RECT 4.400 662.640 1596.000 664.040 ;
        RECT 4.000 650.440 1596.000 662.640 ;
        RECT 4.000 649.040 1595.600 650.440 ;
        RECT 4.000 647.040 1596.000 649.040 ;
        RECT 4.400 645.640 1596.000 647.040 ;
        RECT 4.000 630.040 1596.000 645.640 ;
        RECT 4.000 628.640 1595.600 630.040 ;
        RECT 4.000 626.640 1596.000 628.640 ;
        RECT 4.400 625.240 1596.000 626.640 ;
        RECT 4.000 613.040 1596.000 625.240 ;
        RECT 4.000 611.640 1595.600 613.040 ;
        RECT 4.000 609.640 1596.000 611.640 ;
        RECT 4.400 608.240 1596.000 609.640 ;
        RECT 4.000 596.040 1596.000 608.240 ;
        RECT 4.000 594.640 1595.600 596.040 ;
        RECT 4.000 592.640 1596.000 594.640 ;
        RECT 4.400 591.240 1596.000 592.640 ;
        RECT 4.000 579.040 1596.000 591.240 ;
        RECT 4.000 577.640 1595.600 579.040 ;
        RECT 4.000 575.640 1596.000 577.640 ;
        RECT 4.400 574.240 1596.000 575.640 ;
        RECT 4.000 562.040 1596.000 574.240 ;
        RECT 4.000 560.640 1595.600 562.040 ;
        RECT 4.000 558.640 1596.000 560.640 ;
        RECT 4.400 557.240 1596.000 558.640 ;
        RECT 4.000 545.040 1596.000 557.240 ;
        RECT 4.000 543.640 1595.600 545.040 ;
        RECT 4.000 541.640 1596.000 543.640 ;
        RECT 4.400 540.240 1596.000 541.640 ;
        RECT 4.000 528.040 1596.000 540.240 ;
        RECT 4.000 526.640 1595.600 528.040 ;
        RECT 4.000 524.640 1596.000 526.640 ;
        RECT 4.400 523.240 1596.000 524.640 ;
        RECT 4.000 511.040 1596.000 523.240 ;
        RECT 4.000 509.640 1595.600 511.040 ;
        RECT 4.000 504.240 1596.000 509.640 ;
        RECT 4.400 502.840 1596.000 504.240 ;
        RECT 4.000 490.640 1596.000 502.840 ;
        RECT 4.000 489.240 1595.600 490.640 ;
        RECT 4.000 487.240 1596.000 489.240 ;
        RECT 4.400 485.840 1596.000 487.240 ;
        RECT 4.000 473.640 1596.000 485.840 ;
        RECT 4.000 472.240 1595.600 473.640 ;
        RECT 4.000 470.240 1596.000 472.240 ;
        RECT 4.400 468.840 1596.000 470.240 ;
        RECT 4.000 456.640 1596.000 468.840 ;
        RECT 4.000 455.240 1595.600 456.640 ;
        RECT 4.000 453.240 1596.000 455.240 ;
        RECT 4.400 451.840 1596.000 453.240 ;
        RECT 4.000 439.640 1596.000 451.840 ;
        RECT 4.000 438.240 1595.600 439.640 ;
        RECT 4.000 436.240 1596.000 438.240 ;
        RECT 4.400 434.840 1596.000 436.240 ;
        RECT 4.000 422.640 1596.000 434.840 ;
        RECT 4.000 421.240 1595.600 422.640 ;
        RECT 4.000 419.240 1596.000 421.240 ;
        RECT 4.400 417.840 1596.000 419.240 ;
        RECT 4.000 405.640 1596.000 417.840 ;
        RECT 4.000 404.240 1595.600 405.640 ;
        RECT 4.000 402.240 1596.000 404.240 ;
        RECT 4.400 400.840 1596.000 402.240 ;
        RECT 4.000 388.640 1596.000 400.840 ;
        RECT 4.000 387.240 1595.600 388.640 ;
        RECT 4.000 381.840 1596.000 387.240 ;
        RECT 4.400 380.440 1596.000 381.840 ;
        RECT 4.000 368.240 1596.000 380.440 ;
        RECT 4.000 366.840 1595.600 368.240 ;
        RECT 4.000 364.840 1596.000 366.840 ;
        RECT 4.400 363.440 1596.000 364.840 ;
        RECT 4.000 351.240 1596.000 363.440 ;
        RECT 4.000 349.840 1595.600 351.240 ;
        RECT 4.000 347.840 1596.000 349.840 ;
        RECT 4.400 346.440 1596.000 347.840 ;
        RECT 4.000 334.240 1596.000 346.440 ;
        RECT 4.000 332.840 1595.600 334.240 ;
        RECT 4.000 330.840 1596.000 332.840 ;
        RECT 4.400 329.440 1596.000 330.840 ;
        RECT 4.000 317.240 1596.000 329.440 ;
        RECT 4.000 315.840 1595.600 317.240 ;
        RECT 4.000 313.840 1596.000 315.840 ;
        RECT 4.400 312.440 1596.000 313.840 ;
        RECT 4.000 300.240 1596.000 312.440 ;
        RECT 4.000 298.840 1595.600 300.240 ;
        RECT 4.000 296.840 1596.000 298.840 ;
        RECT 4.400 295.440 1596.000 296.840 ;
        RECT 4.000 283.240 1596.000 295.440 ;
        RECT 4.000 281.840 1595.600 283.240 ;
        RECT 4.000 279.840 1596.000 281.840 ;
        RECT 4.400 278.440 1596.000 279.840 ;
        RECT 4.000 266.240 1596.000 278.440 ;
        RECT 4.000 264.840 1595.600 266.240 ;
        RECT 4.000 262.840 1596.000 264.840 ;
        RECT 4.400 261.440 1596.000 262.840 ;
        RECT 4.000 249.240 1596.000 261.440 ;
        RECT 4.000 247.840 1595.600 249.240 ;
        RECT 4.000 242.440 1596.000 247.840 ;
        RECT 4.400 241.040 1596.000 242.440 ;
        RECT 4.000 228.840 1596.000 241.040 ;
        RECT 4.000 227.440 1595.600 228.840 ;
        RECT 4.000 225.440 1596.000 227.440 ;
        RECT 4.400 224.040 1596.000 225.440 ;
        RECT 4.000 211.840 1596.000 224.040 ;
        RECT 4.000 210.440 1595.600 211.840 ;
        RECT 4.000 208.440 1596.000 210.440 ;
        RECT 4.400 207.040 1596.000 208.440 ;
        RECT 4.000 194.840 1596.000 207.040 ;
        RECT 4.000 193.440 1595.600 194.840 ;
        RECT 4.000 191.440 1596.000 193.440 ;
        RECT 4.400 190.040 1596.000 191.440 ;
        RECT 4.000 177.840 1596.000 190.040 ;
        RECT 4.000 176.440 1595.600 177.840 ;
        RECT 4.000 174.440 1596.000 176.440 ;
        RECT 4.400 173.040 1596.000 174.440 ;
        RECT 4.000 160.840 1596.000 173.040 ;
        RECT 4.000 159.440 1595.600 160.840 ;
        RECT 4.000 157.440 1596.000 159.440 ;
        RECT 4.400 156.040 1596.000 157.440 ;
        RECT 4.000 143.840 1596.000 156.040 ;
        RECT 4.000 142.440 1595.600 143.840 ;
        RECT 4.000 140.440 1596.000 142.440 ;
        RECT 4.400 139.040 1596.000 140.440 ;
        RECT 4.000 126.840 1596.000 139.040 ;
        RECT 4.000 125.440 1595.600 126.840 ;
        RECT 4.000 120.040 1596.000 125.440 ;
        RECT 4.400 118.640 1596.000 120.040 ;
        RECT 4.000 106.440 1596.000 118.640 ;
        RECT 4.000 105.040 1595.600 106.440 ;
        RECT 4.000 103.040 1596.000 105.040 ;
        RECT 4.400 101.640 1596.000 103.040 ;
        RECT 4.000 89.440 1596.000 101.640 ;
        RECT 4.000 88.040 1595.600 89.440 ;
        RECT 4.000 86.040 1596.000 88.040 ;
        RECT 4.400 84.640 1596.000 86.040 ;
        RECT 4.000 72.440 1596.000 84.640 ;
        RECT 4.000 71.040 1595.600 72.440 ;
        RECT 4.000 69.040 1596.000 71.040 ;
        RECT 4.400 67.640 1596.000 69.040 ;
        RECT 4.000 55.440 1596.000 67.640 ;
        RECT 4.000 54.040 1595.600 55.440 ;
        RECT 4.000 52.040 1596.000 54.040 ;
        RECT 4.400 50.640 1596.000 52.040 ;
        RECT 4.000 38.440 1596.000 50.640 ;
        RECT 4.000 37.040 1595.600 38.440 ;
        RECT 4.000 35.040 1596.000 37.040 ;
        RECT 4.400 33.640 1596.000 35.040 ;
        RECT 4.000 21.440 1596.000 33.640 ;
        RECT 4.000 20.040 1595.600 21.440 ;
        RECT 4.000 18.040 1596.000 20.040 ;
        RECT 4.400 16.640 1596.000 18.040 ;
        RECT 4.000 4.440 1596.000 16.640 ;
        RECT 4.000 3.575 1595.600 4.440 ;
      LAYER met4 ;
        RECT 279.975 19.895 327.840 1587.625 ;
        RECT 330.240 19.895 404.640 1587.625 ;
        RECT 407.040 19.895 481.440 1587.625 ;
        RECT 483.840 19.895 558.240 1587.625 ;
        RECT 560.640 19.895 635.040 1587.625 ;
        RECT 637.440 19.895 711.840 1587.625 ;
        RECT 714.240 19.895 788.640 1587.625 ;
        RECT 791.040 19.895 865.440 1587.625 ;
        RECT 867.840 19.895 942.240 1587.625 ;
        RECT 944.640 19.895 1019.040 1587.625 ;
        RECT 1021.440 19.895 1095.840 1587.625 ;
        RECT 1098.240 19.895 1172.640 1587.625 ;
        RECT 1175.040 19.895 1249.440 1587.625 ;
        RECT 1251.840 19.895 1326.240 1587.625 ;
        RECT 1328.640 19.895 1403.040 1587.625 ;
        RECT 1405.440 19.895 1479.840 1587.625 ;
        RECT 1482.240 19.895 1556.640 1587.625 ;
        RECT 1559.040 19.895 1577.505 1587.625 ;
  END
END core_empty
END LIBRARY

